VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO scs130lp_a2111o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111o_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.915 0.78 3.25 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.42 0.78 3.755 1.845 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.04 1.135 2.41 2.27 ;
        RECT 2.04 1.135 2.245 2.54 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.135 1.87 2.94 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.98 1.135 1.375 1.875 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.28 0.645 0.61 ;
        RECT 0.085 0.28 0.365 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.215 -0.085 3.595 0.61 ;
        RECT 1.68 -0.085 2.32 0.61 ;
        RECT 0.815 -0.085 1.075 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.99 2.37 3.255 3.415 ;
        RECT 0.535 2.405 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.425 2.02 3.72 3.04 ;
      RECT 2.315 2.71 2.82 3.04 ;
      RECT 2.58 2.02 2.82 3.04 ;
      RECT 2.58 2.02 3.72 2.19 ;
      RECT 1.105 2.055 1.375 3.04 ;
      RECT 0.535 2.055 1.375 2.225 ;
      RECT 0.535 0.795 0.81 2.225 ;
      RECT 0.535 0.795 2.745 0.965 ;
      RECT 2.49 0.28 2.745 0.965 ;
      RECT 1.245 0.28 1.51 0.965 ;
  END
END scs130lp_a2111o_0

MACRO scs130lp_a2111o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111o_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.99 1.21 3.695 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.865 1.21 4.235 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.435 1.335 2.82 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 1.335 2.265 2.96 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.075 1.335 1.775 1.75 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.255 0.52 1.775 ;
        RECT 0.085 0.255 0.48 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.7 -0.085 4.03 1.04 ;
        RECT 2.03 -0.085 2.36 0.825 ;
        RECT 0.69 -0.085 1.46 0.825 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.3 2.27 3.63 3.415 ;
        RECT 0.65 2.26 0.98 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.8 1.93 4.06 3.075 ;
      RECT 2.53 1.93 3.13 3.075 ;
      RECT 2.53 1.93 4.06 2.1 ;
      RECT 1.17 1.92 1.5 3.075 ;
      RECT 0.69 1.92 1.5 2.09 ;
      RECT 0.69 0.995 0.905 2.09 ;
      RECT 0.69 0.995 2.82 1.165 ;
      RECT 2.53 0.255 3.24 1.04 ;
      RECT 1.63 0.255 1.86 1.165 ;
  END
END scs130lp_a2111o_1

MACRO scs130lp_a2111o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111o_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 0.3 3.775 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.945 1.21 4.715 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.965 1.345 3.31 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.345 2.795 2.965 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.345 2.255 1.75 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.255 0.895 2.1 ;
        RECT 0.625 0.255 0.815 3 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.09 -0.085 4.42 1.04 ;
        RECT 2.59 -0.085 2.92 0.815 ;
        RECT 1.065 -0.085 2.01 0.835 ;
        RECT 0.205 -0.085 0.455 1.105 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.605 2.27 3.935 3.415 ;
        RECT 0.985 2.27 1.315 3.415 ;
        RECT 0.125 1.815 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.105 1.93 4.42 3.075 ;
      RECT 3.07 1.93 3.4 3.075 ;
      RECT 3.07 1.93 4.42 2.1 ;
      RECT 1.68 1.92 2.01 3.075 ;
      RECT 1.065 1.92 2.01 2.1 ;
      RECT 1.065 1.005 1.415 2.1 ;
      RECT 1.065 1.005 3.335 1.175 ;
      RECT 3.09 0.255 3.335 1.175 ;
      RECT 2.18 0.255 2.42 1.175 ;
  END
END scs130lp_a2111o_2

MACRO scs130lp_a2111o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111o_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.695 1.21 5.17 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.34 1.21 5.85 1.445 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.375 1.335 4.165 1.785 ;
        RECT 2.965 1.335 4.165 1.535 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.425 2.795 1.77 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.425 0.535 1.75 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.39 1.745 8.075 1.925 ;
        RECT 7.715 1.065 8.075 1.925 ;
        RECT 6.39 1.065 8.075 1.235 ;
        RECT 7.25 1.745 7.44 3.075 ;
        RECT 7.25 0.255 7.44 1.235 ;
        RECT 6.39 1.745 6.58 3.075 ;
        RECT 6.39 0.255 6.58 1.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.61 -0.085 7.94 0.895 ;
        RECT 6.75 -0.085 7.08 0.895 ;
        RECT 5.89 -0.085 6.22 1.04 ;
        RECT 5.03 -0.085 5.36 0.59 ;
        RECT 2.575 -0.085 3.51 0.815 ;
        RECT 1.675 -0.085 2.005 0.815 ;
        RECT 0.775 -0.085 1.105 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.61 2.105 7.94 3.415 ;
        RECT 6.75 2.095 7.08 3.415 ;
        RECT 5.89 1.955 6.22 3.415 ;
        RECT 5.03 2.295 5.36 3.415 ;
        RECT 4.04 2.295 4.37 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.705 1.93 1.035 2.735 ;
      RECT 0.705 1.065 0.935 2.735 ;
      RECT 4.345 1.615 6.2 1.785 ;
      RECT 6.02 1.405 6.2 1.785 ;
      RECT 4.345 0.985 4.515 1.785 ;
      RECT 6.02 1.405 7.545 1.575 ;
      RECT 0.345 1.065 1.455 1.235 ;
      RECT 1.275 0.985 4.515 1.155 ;
      RECT 0.345 0.255 0.605 1.235 ;
      RECT 3.68 0.255 3.87 1.155 ;
      RECT 2.175 0.255 2.405 1.155 ;
      RECT 1.275 0.255 1.505 1.155 ;
      RECT 3.68 0.255 4.8 0.465 ;
      RECT 4.685 0.76 5.72 1.04 ;
      RECT 5.53 0.255 5.72 1.04 ;
      RECT 4.04 0.635 4.86 0.815 ;
      RECT 5.53 1.955 5.72 3.075 ;
      RECT 2.515 2.905 3.825 3.075 ;
      RECT 3.495 1.955 3.825 3.075 ;
      RECT 4.54 1.955 4.8 3.025 ;
      RECT 2.515 2.28 2.845 3.075 ;
      RECT 3.495 1.955 5.72 2.125 ;
      RECT 3.015 1.705 3.205 2.735 ;
      RECT 1.565 1.94 1.895 2.735 ;
      RECT 1.565 1.94 3.205 2.11 ;
      RECT 2.965 1.705 3.205 2.11 ;
      RECT 0.275 2.905 2.325 3.075 ;
      RECT 2.065 2.28 2.325 3.075 ;
      RECT 1.205 1.94 1.395 3.075 ;
      RECT 0.275 1.92 0.535 3.075 ;
  END
END scs130lp_a2111o_4

MACRO scs130lp_a2111o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111o_lp 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 1.175 5.155 1.845 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.935 1.175 4.265 1.845 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.365 1.175 3.715 1.845 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 1.175 1.39 1.845 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.855 0.53 1.78 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.235 0.265 2.845 0.645 ;
        RECT 2.235 1.92 2.755 2.18 ;
        RECT 2.235 0.265 2.405 2.18 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 3.885 -0.085 4.215 0.645 ;
        RECT 1.725 -0.085 2.055 0.645 ;
        RECT 0.115 -0.085 0.445 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.2 2.375 4.53 3.415 ;
        RECT 1.835 2.71 2.165 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.805 2.025 5.135 3.065 ;
      RECT 3.67 2.025 4 3.065 ;
      RECT 3.67 2.025 5.135 2.195 ;
      RECT 2.585 0.825 2.915 1.495 ;
      RECT 2.585 0.825 5.035 0.995 ;
      RECT 4.705 0.265 5.035 0.995 ;
      RECT 3.095 0.265 3.425 0.995 ;
      RECT 3.14 2.025 3.47 3.065 ;
      RECT 1.135 2.025 1.465 3.065 ;
      RECT 1.135 2.36 3.47 2.53 ;
      RECT 0.115 2.025 0.445 3.065 ;
      RECT 0.115 2.025 0.88 2.195 ;
      RECT 0.71 0.265 0.88 2.195 ;
      RECT 1.725 0.825 2.055 1.79 ;
      RECT 0.71 0.825 2.055 0.995 ;
      RECT 0.71 0.265 1.265 0.995 ;
  END
END scs130lp_a2111o_lp

MACRO scs130lp_a2111o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111o_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.7 2.665 3.205 2.995 ;
        RECT 2.89 2.32 3.205 2.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.84 3.205 1.38 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 2.735 2.17 3.065 ;
        RECT 1.5 2.32 1.765 3.065 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 2.32 1.33 2.965 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.965 1.095 1.295 1.75 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.53 0.39 2.86 ;
        RECT 0.155 0.345 0.39 0.675 ;
        RECT 0.155 0.345 0.325 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.85 -0.085 3.18 0.485 ;
        RECT 1.69 -0.085 1.9 0.545 ;
        RECT 0.57 -0.085 0.9 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.52 1.955 2.71 2.495 ;
        RECT 2.34 2.305 2.53 3.415 ;
        RECT 0.61 2.645 0.82 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.09 1.605 2.3 2.135 ;
      RECT 2.93 1.605 3.26 2.095 ;
      RECT 2.09 1.605 3.26 1.775 ;
      RECT 0.505 1.93 1.645 2.14 ;
      RECT 1.475 0.725 1.645 2.14 ;
      RECT 0.505 1.47 0.675 2.14 ;
      RECT 1.26 0.725 2.33 0.895 ;
      RECT 2.12 0.345 2.33 0.895 ;
      RECT 1.26 0.345 1.47 0.895 ;
  END
END scs130lp_a2111o_m

MACRO scs130lp_a2111oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111oi_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.435 0.78 2.765 1.875 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 0.84 3.275 2.225 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.19 2.265 1.86 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.98 1.19 1.35 2.93 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.365 2.21 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.535 0.78 2.265 1.02 ;
        RECT 1.735 0.28 2.265 1.02 ;
        RECT 0.81 0.28 1.065 1.02 ;
        RECT 0.385 2.395 0.705 3.065 ;
        RECT 0.535 0.78 0.705 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.495 -0.085 2.825 0.61 ;
        RECT 1.235 -0.085 1.56 0.61 ;
        RECT 0.345 -0.085 0.64 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.04 2.405 2.37 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.54 2.395 2.855 3.065 ;
      RECT 1.565 2.045 1.86 3.065 ;
      RECT 2.54 2.045 2.765 3.065 ;
      RECT 1.565 2.045 2.765 2.225 ;
  END
END scs130lp_a2111oi_0

MACRO scs130lp_a2111oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111oi_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.185 2.725 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.19 3.27 1.52 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.485 1.185 1.875 1.52 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.21 1.315 3.02 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.535 1.345 0.855 2.86 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2894 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.97 0.255 2.725 1.015 ;
        RECT 0.635 0.84 2.725 1.015 ;
        RECT 0.635 0.255 0.965 1.015 ;
        RECT 0.115 0.985 0.855 1.155 ;
        RECT 0.115 0.985 0.365 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.895 -0.085 3.16 1.015 ;
        RECT 1.135 -0.085 1.8 0.67 ;
        RECT 0.135 -0.085 0.465 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.325 2.105 2.655 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.89 1.755 3.16 3.075 ;
      RECT 1.765 1.755 2.095 3.075 ;
      RECT 1.765 1.755 3.16 1.925 ;
  END
END scs130lp_a2111oi_1

MACRO scs130lp_a2111oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111oi_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.465 1.615 5.155 1.785 ;
        RECT 4.895 1.345 5.155 1.785 ;
        RECT 3.465 1.345 4.185 1.785 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.355 1.21 4.725 1.435 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.425 2.855 1.775 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.605 1.895 1.775 ;
        RECT 1.525 1.295 1.895 1.775 ;
        RECT 0.125 1.295 0.455 1.775 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.21 1.355 1.435 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5414 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 1.955 5.66 2.125 ;
        RECT 5.325 0.255 5.66 2.125 ;
        RECT 5.02 0.255 5.66 1.095 ;
        RECT 1 1.945 3.295 2.125 ;
        RECT 3.025 0.255 3.295 2.125 ;
        RECT 2.065 1.085 3.295 1.255 ;
        RECT 2.965 0.255 3.295 1.255 ;
        RECT 2.065 0.255 2.295 1.255 ;
        RECT 0.12 0.87 2.295 1.04 ;
        RECT 1.965 0.255 2.295 1.04 ;
        RECT 1.05 0.265 1.295 1.04 ;
        RECT 1 1.945 1.265 2.355 ;
        RECT 0.12 0.255 0.38 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.125 -0.085 4.455 0.7 ;
        RECT 2.465 -0.085 2.795 0.915 ;
        RECT 1.465 -0.085 1.795 0.7 ;
        RECT 0.55 -0.085 0.88 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.57 2.635 4.9 3.415 ;
        RECT 3.69 2.635 4.02 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.07 2.295 5.35 3.075 ;
      RECT 4.19 2.295 4.4 3.075 ;
      RECT 3.26 2.295 3.52 3.075 ;
      RECT 2.335 2.295 3.52 2.645 ;
      RECT 2.335 2.295 5.35 2.465 ;
      RECT 3.53 0.87 4.85 1.04 ;
      RECT 4.625 0.255 4.85 1.04 ;
      RECT 3.53 0.255 3.86 1.04 ;
      RECT 0.12 2.865 3.07 3.075 ;
      RECT 1.87 2.815 3.07 3.075 ;
      RECT 0.12 1.955 0.4 3.075 ;
      RECT 1.87 2.295 2.165 3.075 ;
      RECT 0.57 2.525 1.7 2.695 ;
      RECT 1.45 2.295 1.7 2.695 ;
      RECT 0.57 1.955 0.83 2.695 ;
  END
END scs130lp_a2111oi_2

MACRO scs130lp_a2111oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111oi_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.845 1.21 7.7 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.945 1.375 9.975 1.545 ;
        RECT 7.945 1.375 8.485 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.95 1.425 5.675 1.76 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.05 1.425 3.74 1.76 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.49 1.21 1.84 1.435 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.945 0.87 7.605 1.04 ;
        RECT 7.31 0.595 7.605 1.04 ;
        RECT 6.46 0.595 6.705 1.04 ;
        RECT 4.945 0.255 5.195 1.04 ;
        RECT 2.305 1.085 5.185 1.255 ;
        RECT 4.945 0.255 5.185 1.255 ;
        RECT 4.095 0.255 4.335 1.255 ;
        RECT 3.175 0.255 3.425 1.255 ;
        RECT 2.305 0.87 2.505 1.255 ;
        RECT 2.315 0.255 2.505 1.255 ;
        RECT 0.14 0.87 2.505 1.04 ;
        RECT 1.455 1.705 1.645 2.735 ;
        RECT 1.455 0.255 1.645 1.04 ;
        RECT 0.14 1.705 1.645 1.875 ;
        RECT 0.595 1.705 0.785 2.735 ;
        RECT 0.595 0.255 0.785 1.04 ;
        RECT 0.14 0.87 0.32 1.875 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.09 -0.085 9.42 0.865 ;
        RECT 8.23 -0.085 8.56 0.865 ;
        RECT 5.365 -0.085 5.695 0.69 ;
        RECT 4.505 -0.085 4.775 0.915 ;
        RECT 3.595 -0.085 3.925 0.915 ;
        RECT 2.675 -0.085 3.005 0.915 ;
        RECT 1.815 -0.085 2.145 0.7 ;
        RECT 0.955 -0.085 1.285 0.7 ;
        RECT 0.095 -0.085 0.425 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.015 2.055 9.345 3.415 ;
        RECT 8.065 2.27 8.395 3.415 ;
        RECT 7.065 1.945 7.395 3.415 ;
        RECT 6.205 1.945 6.535 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 7.87 1.035 9.85 1.205 ;
      RECT 9.59 0.255 9.85 1.205 ;
      RECT 8.73 0.255 8.92 1.205 ;
      RECT 7.87 0.255 8.06 1.205 ;
      RECT 6.875 0.255 7.14 0.7 ;
      RECT 5.965 0.255 6.29 0.7 ;
      RECT 5.965 0.255 8.06 0.425 ;
      RECT 9.515 1.715 9.775 3.075 ;
      RECT 8.565 1.93 8.845 3.075 ;
      RECT 8.655 1.715 8.845 3.075 ;
      RECT 7.565 1.93 7.895 3.075 ;
      RECT 6.705 1.605 6.895 3.075 ;
      RECT 4.055 2.905 6.035 3.075 ;
      RECT 5.845 1.605 6.035 3.075 ;
      RECT 4.955 2.305 5.175 3.075 ;
      RECT 4.055 2.27 4.385 3.075 ;
      RECT 7.565 1.93 8.845 2.1 ;
      RECT 7.565 1.605 7.775 3.075 ;
      RECT 8.655 1.715 9.775 1.885 ;
      RECT 5.845 1.605 7.775 1.775 ;
      RECT 5.345 1.93 5.675 2.735 ;
      RECT 4.555 1.93 4.785 2.735 ;
      RECT 3.175 1.93 3.365 2.735 ;
      RECT 2.315 1.93 2.505 2.735 ;
      RECT 4.555 1.93 5.675 2.12 ;
      RECT 2.315 1.93 5.675 2.1 ;
      RECT 0.095 2.905 3.865 3.075 ;
      RECT 3.535 2.27 3.865 3.075 ;
      RECT 2.675 2.27 3.005 3.075 ;
      RECT 1.815 1.93 2.145 3.075 ;
      RECT 0.955 2.045 1.285 3.075 ;
      RECT 0.095 2.045 0.425 3.075 ;
  END
END scs130lp_a2111oi_4

MACRO scs130lp_a2111oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111oi_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.175 0.835 1.845 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.175 1.795 1.845 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.175 2.755 1.845 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 1.18 3.265 2.89 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 1.175 3.835 1.845 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6357 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.73 2.025 4.185 3.065 ;
        RECT 4.015 0.825 4.185 3.065 ;
        RECT 0.17 0.825 4.185 0.995 ;
        RECT 3.005 0.265 3.43 0.995 ;
        RECT 1.78 0.265 2.11 0.995 ;
        RECT 0.17 0.265 0.5 0.995 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.89 -0.085 4.22 0.645 ;
        RECT 2.31 -0.085 2.64 0.645 ;
        RECT 0.99 -0.085 1.32 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 1.16 2.375 1.49 3.415 ;
        RECT 0.1 2.025 0.43 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.14 2.025 2.47 3.065 ;
      RECT 0.63 2.025 0.96 3.065 ;
      RECT 0.63 2.025 2.47 2.195 ;
  END
END scs130lp_a2111oi_lp

MACRO scs130lp_a2111oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2111oi_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.315 2.195 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3 0.47 3.205 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.775 2.12 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.975 1.315 2.12 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 1.21 0.805 2.86 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.441 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.82 0.345 2.03 0.795 ;
        RECT 0.635 0.625 2.03 0.795 ;
        RECT 0.635 0.345 1.02 0.795 ;
        RECT 0.155 0.725 0.805 0.895 ;
        RECT 0.155 0.725 0.345 2.975 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.61 -0.085 2.82 0.545 ;
        RECT 1.2 -0.085 1.53 0.445 ;
        RECT 0.265 -0.085 0.455 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.92 2.835 2.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.53 2.485 1.74 2.975 ;
      RECT 2.55 2.485 2.88 2.915 ;
      RECT 1.53 2.485 2.88 2.655 ;
  END
END scs130lp_a2111oi_m

MACRO scs130lp_a211o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211o_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.2 1.835 1.89 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 1.2 1.345 1.88 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.2 2.365 1.88 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.875 1.2 3.275 2.195 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 0.345 0.39 0.675 ;
        RECT 0.095 2.18 0.385 2.935 ;
        RECT 0.095 0.345 0.335 2.935 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.13 -0.085 2.72 0.675 ;
        RECT 0.56 -0.085 1.2 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.55 2.4 1.84 3.415 ;
        RECT 0.555 2.18 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.615 2.39 3.1 3.06 ;
      RECT 2.535 0.86 2.705 2.56 ;
      RECT 0.505 0.86 0.755 1.53 ;
      RECT 0.505 0.86 3.19 1.03 ;
      RECT 2.89 0.345 3.19 1.03 ;
      RECT 1.66 0.345 1.96 1.03 ;
      RECT 2.01 2.06 2.275 3.075 ;
      RECT 1.08 2.06 1.38 3.07 ;
      RECT 1.08 2.06 2.275 2.23 ;
  END
END scs130lp_a211o_0

MACRO scs130lp_a211o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211o_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.21 2.04 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.195 1.39 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.25 1.21 2.735 1.525 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.21 3.235 1.525 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 0.255 0.405 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.445 -0.085 2.775 0.685 ;
        RECT 0.575 -0.085 1.345 0.685 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.515 2.375 1.845 3.415 ;
        RECT 0.575 2.045 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.915 1.695 3.245 3.075 ;
      RECT 0.585 1.695 3.245 1.865 ;
      RECT 0.585 0.855 0.915 1.865 ;
      RECT 0.585 0.855 3.245 1.025 ;
      RECT 2.945 0.255 3.245 1.025 ;
      RECT 1.905 0.255 2.235 1.025 ;
      RECT 2.03 2.035 2.36 3.075 ;
      RECT 1.045 2.035 1.345 3.075 ;
      RECT 1.045 2.035 2.36 2.205 ;
  END
END scs130lp_a211o_1

MACRO scs130lp_a211o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211o_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 1.195 2.47 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.195 1.845 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.68 1.195 3.215 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.195 3.755 1.515 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 0.255 0.825 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.915 -0.085 3.245 0.685 ;
        RECT 0.995 -0.085 1.805 0.685 ;
        RECT 0.095 -0.085 0.385 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.96 2.395 2.29 3.415 ;
        RECT 1 2.045 1.285 3.415 ;
        RECT 0.095 1.815 0.385 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.345 1.695 3.675 3.075 ;
      RECT 1.245 1.695 3.675 1.875 ;
      RECT 1.245 0.855 1.415 1.875 ;
      RECT 1 1.345 1.415 1.675 ;
      RECT 1.245 0.855 3.675 1.025 ;
      RECT 3.415 0.255 3.675 1.025 ;
      RECT 2.365 0.255 2.695 1.025 ;
      RECT 1.475 2.045 1.79 3.075 ;
      RECT 2.46 2.045 2.79 3.065 ;
      RECT 1.475 2.045 2.79 2.225 ;
  END
END scs130lp_a211o_2

MACRO scs130lp_a211o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211o_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.31 1.425 5.64 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.915 1.345 6.5 1.645 ;
        RECT 4.9 1.95 6.125 2.12 ;
        RECT 5.915 1.345 6.125 2.12 ;
        RECT 4.9 1.425 5.1 2.12 ;
        RECT 4.77 1.425 5.1 1.82 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.815 1.695 4.45 1.865 ;
        RECT 4.12 1.415 4.45 1.865 ;
        RECT 2.815 1.345 3.205 1.865 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.375 1.185 3.71 1.515 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1886 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 1.055 2.305 1.225 ;
        RECT 2.125 0.255 2.305 1.225 ;
        RECT 1.265 1.045 2.305 1.225 ;
        RECT 1.57 1.755 1.76 3.075 ;
        RECT 0.09 1.755 1.76 1.925 ;
        RECT 1.265 0.255 1.455 1.225 ;
        RECT 0.71 1.755 0.9 3.075 ;
        RECT 0.09 0.39 0.405 1.225 ;
        RECT 0.09 0.39 0.345 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 6.365 -0.085 6.625 1.095 ;
        RECT 4.28 -0.085 4.835 0.885 ;
        RECT 3.375 -0.085 3.705 0.675 ;
        RECT 2.5 -0.085 2.83 0.805 ;
        RECT 1.625 -0.085 1.955 0.875 ;
        RECT 0.765 -0.085 1.095 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.865 2.63 6.195 3.415 ;
        RECT 4.895 2.63 5.225 3.415 ;
        RECT 1.93 1.815 2.26 3.415 ;
        RECT 1.07 2.105 1.4 3.415 ;
        RECT 0.21 2.095 0.54 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.365 1.815 6.625 3.075 ;
      RECT 5.435 2.29 5.695 3.075 ;
      RECT 4.385 2.035 4.725 3.075 ;
      RECT 2.595 2.375 2.855 3.075 ;
      RECT 2.595 2.425 4.725 2.595 ;
      RECT 6.295 1.815 6.625 2.46 ;
      RECT 4.355 2.29 6.625 2.46 ;
      RECT 2.595 2.375 2.925 2.595 ;
      RECT 4.355 2.035 4.73 2.46 ;
      RECT 5.865 0.255 6.195 1.095 ;
      RECT 5.005 0.255 5.335 0.895 ;
      RECT 5.005 0.255 6.195 0.425 ;
      RECT 3.455 2.035 3.785 2.255 ;
      RECT 2.475 2.035 3.785 2.205 ;
      RECT 2.475 0.985 2.645 2.205 ;
      RECT 0.515 1.395 2.645 1.585 ;
      RECT 3.885 1.065 5.695 1.235 ;
      RECT 5.505 0.595 5.695 1.235 ;
      RECT 2.475 0.985 3.205 1.155 ;
      RECT 3 0.255 3.205 1.155 ;
      RECT 3.885 0.255 4.11 1.235 ;
      RECT 3.875 0.255 4.11 1.015 ;
      RECT 3 0.845 4.11 1.015 ;
      RECT 3.025 2.765 4.215 3.055 ;
  END
END scs130lp_a211o_4

MACRO scs130lp_a211o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211o_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.955 0.485 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.93 1.17 1.315 1.84 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 1.17 1.83 1.84 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.17 2.4 1.84 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 0.265 3.715 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.595 -0.085 2.925 0.64 ;
        RECT 1.015 -0.085 1.345 0.64 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.855 2.37 3.185 3.415 ;
        RECT 0.655 2.37 0.985 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.295 2.02 2.625 3.065 ;
      RECT 2.295 2.02 3.045 2.19 ;
      RECT 2.875 0.82 3.045 2.19 ;
      RECT 2.875 0.82 3.205 1.49 ;
      RECT 0.665 0.82 3.205 0.99 ;
      RECT 1.805 0.265 2.135 0.99 ;
      RECT 0.665 0.555 0.835 0.99 ;
      RECT 0.195 0.555 0.835 0.725 ;
      RECT 0.195 0.265 0.525 0.725 ;
      RECT 1.235 2.02 1.565 3.065 ;
      RECT 0.125 2.02 0.455 3.065 ;
      RECT 0.125 2.02 1.565 2.19 ;
  END
END scs130lp_a211o_lp

MACRO scs130lp_a211o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211o_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.265 1.285 1.01 ;
        RECT 0.92 0.265 1.285 0.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.33 1.21 1.765 1.585 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.265 2.43 0.595 ;
        RECT 1.595 0.265 2.245 0.64 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.76 1.535 3.205 1.75 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.47 0.39 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.455 0.775 2.785 0.985 ;
        RECT 2.615 -0.085 2.785 0.985 ;
        RECT 0.57 0.765 0.9 0.975 ;
        RECT 0.57 -0.085 0.74 0.975 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.515 2.115 1.845 3.415 ;
        RECT 0.595 2.785 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.025 2.735 2.565 3.065 ;
      RECT 2.395 1.165 2.565 3.065 ;
      RECT 2.395 1.93 3.005 2.26 ;
      RECT 1.945 1.165 3.155 1.335 ;
      RECT 2.965 0.835 3.155 1.335 ;
      RECT 1.945 0.915 2.275 1.335 ;
      RECT 2.025 1.765 2.215 2.255 ;
      RECT 1.145 1.765 1.335 2.255 ;
      RECT 1.145 1.765 2.215 1.935 ;
  END
END scs130lp_a211o_m

MACRO scs130lp_a211oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211oi_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 0.78 0.98 1.875 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.425 1.875 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.47 1.155 1.815 1.825 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.385 1.21 2.795 2.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5413 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 0.28 2.795 1.04 ;
        RECT 1.925 2.395 2.215 3.075 ;
        RECT 1.985 0.78 2.215 3.075 ;
        RECT 1.15 0.78 2.795 0.985 ;
        RECT 1.15 0.28 1.4 0.985 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.57 -0.085 1.83 0.61 ;
        RECT 0.285 -0.085 0.615 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 0.71 2.395 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.14 2.045 1.435 3.075 ;
      RECT 0.245 2.045 0.54 3.075 ;
      RECT 0.245 2.045 1.435 2.225 ;
  END
END scs130lp_a211oi_0

MACRO scs130lp_a211oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211oi_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.195 1.01 1.525 ;
        RECT 0.595 1.195 0.875 1.76 ;
        RECT 0.595 0.38 0.845 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.21 0.425 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.265 1.345 1.8 1.76 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.97 1.345 2.305 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8841 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.965 1.925 2.785 3.075 ;
        RECT 2.5 0.885 2.785 3.075 ;
        RECT 1.18 0.995 2.785 1.175 ;
        RECT 2.02 0.885 2.785 1.175 ;
        RECT 2.02 0.255 2.295 1.175 ;
        RECT 1.18 0.255 1.35 1.175 ;
        RECT 1.015 0.255 1.35 0.965 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.52 -0.085 1.85 0.825 ;
        RECT 0.095 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 0.58 2.27 0.91 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.125 1.93 1.455 3.075 ;
      RECT 0.095 1.93 0.41 3.075 ;
      RECT 0.095 1.93 1.455 2.1 ;
  END
END scs130lp_a211oi_1

MACRO scs130lp_a211oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211oi_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 1.21 4.715 1.75 ;
        RECT 3.73 1.415 4.715 1.595 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.415 3.45 1.595 ;
        RECT 2.005 1.415 2.895 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.425 1.835 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.425 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1256 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.075 4.265 1.245 ;
        RECT 3.935 0.595 4.265 1.245 ;
        RECT 1.525 0.255 1.765 1.245 ;
        RECT 0.595 1.075 0.925 2.735 ;
        RECT 0.595 0.255 0.855 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 2.915 -0.085 3.245 0.565 ;
        RECT 1.935 -0.085 2.215 0.905 ;
        RECT 1.025 -0.085 1.355 0.905 ;
        RECT 0.165 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.285 1.92 4.615 3.415 ;
        RECT 3.425 2.105 3.755 3.415 ;
        RECT 2.565 2.26 2.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.435 0.255 4.695 1.04 ;
      RECT 2.405 0.735 3.755 0.905 ;
      RECT 3.425 0.255 3.755 0.905 ;
      RECT 2.405 0.305 2.735 0.905 ;
      RECT 3.425 0.255 4.695 0.425 ;
      RECT 3.925 1.765 4.115 3.075 ;
      RECT 3.065 1.765 3.255 3.075 ;
      RECT 1.455 1.92 1.785 2.735 ;
      RECT 1.455 1.92 3.255 2.09 ;
      RECT 3.065 1.765 4.115 1.935 ;
      RECT 0.165 2.905 2.215 3.075 ;
      RECT 1.955 2.26 2.215 3.075 ;
      RECT 1.095 1.92 1.285 3.075 ;
      RECT 0.165 1.92 0.425 3.075 ;
  END
END scs130lp_a211oi_2

MACRO scs130lp_a211oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211oi_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.835 1.18 3.205 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.27 3.76 1.535 ;
        RECT 0.12 1.615 3.555 1.785 ;
        RECT 3.385 1.27 3.555 1.785 ;
        RECT 0.12 1.345 1.645 1.785 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.98 1.085 7.24 1.515 ;
        RECT 4.895 1.085 7.24 1.255 ;
        RECT 3.98 1.21 5.18 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.35 1.425 6.71 1.645 ;
        RECT 5.35 1.425 6.145 1.765 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.1168 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.41 0.745 7.58 1.985 ;
        RECT 6.315 1.815 7.58 1.985 ;
        RECT 4.055 0.745 7.58 0.915 ;
        RECT 6.675 0.255 7.005 0.915 ;
        RECT 5.395 1.935 6.615 2.145 ;
        RECT 5.815 0.255 6.145 0.915 ;
        RECT 4.055 0.725 5.285 0.915 ;
        RECT 4.955 0.255 5.285 0.915 ;
        RECT 1.835 0.755 4.725 1.01 ;
        RECT 4.055 0.255 4.355 1.01 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.175 -0.085 7.435 0.575 ;
        RECT 6.315 -0.085 6.505 0.575 ;
        RECT 5.455 -0.085 5.645 0.575 ;
        RECT 4.525 -0.085 4.785 0.555 ;
        RECT 3.555 -0.085 3.885 0.585 ;
        RECT 0.975 -0.085 1.305 0.835 ;
        RECT 0.115 -0.085 0.415 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 3.195 2.295 3.525 3.415 ;
        RECT 2.335 2.295 2.665 3.415 ;
        RECT 1.475 2.295 1.805 3.415 ;
        RECT 0.615 2.295 0.945 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.695 1.955 3.945 3.075 ;
      RECT 3.735 1.705 3.945 3.075 ;
      RECT 2.835 1.955 3.025 3.075 ;
      RECT 1.975 1.955 2.165 3.075 ;
      RECT 1.115 1.955 1.305 3.075 ;
      RECT 0.185 1.955 0.445 3.075 ;
      RECT 7.135 2.165 7.465 3.055 ;
      RECT 4.595 2.325 7.465 2.575 ;
      RECT 4.595 1.705 4.805 2.575 ;
      RECT 0.185 1.955 3.945 2.125 ;
      RECT 3.735 1.705 4.805 1.875 ;
      RECT 4.165 2.745 6.965 3.075 ;
      RECT 4.165 2.045 4.375 3.075 ;
      RECT 0.585 1.005 1.665 1.175 ;
      RECT 1.475 0.255 1.665 1.175 ;
      RECT 0.585 0.255 0.805 1.175 ;
      RECT 1.475 0.255 3.385 0.585 ;
  END
END scs130lp_a211oi_4

MACRO scs130lp_a211oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211oi_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.17 2.305 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.11 3.235 1.78 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.17 1.795 1.84 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 1.18 0.905 2.89 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7273 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.82 2.14 0.99 ;
        RECT 1.81 0.265 2.14 0.99 ;
        RECT 0.125 0.265 0.56 0.99 ;
        RECT 0.125 0.265 0.395 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.67 -0.085 3 0.725 ;
        RECT 1.02 -0.085 1.35 0.64 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.94 2.37 2.27 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.77 2.02 3.1 3.065 ;
      RECT 1.41 2.02 1.74 3.065 ;
      RECT 1.41 2.02 3.1 2.19 ;
  END
END scs130lp_a211oi_lp

MACRO scs130lp_a211oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a211oi_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.995 1.09 1.505 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.84 0.455 1.38 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.3 0.995 1.765 1.505 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.32 2.605 2.245 2.945 ;
        RECT 1.85 2.32 2.245 2.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3864 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.965 0.645 2.295 2.12 ;
        RECT 2.025 0.345 2.295 2.12 ;
        RECT 1.055 0.645 2.295 0.815 ;
        RECT 1.055 0.345 1.265 0.815 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.445 -0.085 1.775 0.465 ;
        RECT 0.095 -0.085 0.425 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.545 2.035 0.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.155 1.685 0.365 2.155 ;
      RECT 1.125 1.685 1.335 2.135 ;
      RECT 0.155 1.685 1.335 1.855 ;
  END
END scs130lp_a211oi_m

MACRO scs130lp_a21bo_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21bo_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 0.805 2.795 1.755 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.965 0.805 3.375 1.76 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.93 0.83 1.33 1.39 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 0.305 0.535 0.635 ;
        RECT 0.09 1.95 0.42 3.06 ;
        RECT 0.09 0.305 0.26 3.06 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.17 -0.085 3.5 0.635 ;
        RECT 1.84 -0.085 2.035 0.635 ;
        RECT 0.705 -0.085 0.955 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.77 2.28 3.035 3.415 ;
        RECT 0.59 2.4 0.885 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.205 1.93 3.5 2.94 ;
      RECT 2.34 1.93 2.6 2.94 ;
      RECT 2.34 1.93 3.5 2.1 ;
      RECT 1.88 1.56 2.17 2.94 ;
      RECT 0.43 1.56 2.375 1.73 ;
      RECT 2.205 0.305 2.375 1.73 ;
      RECT 0.43 1.06 0.695 1.73 ;
      RECT 2.205 0.305 2.54 0.635 ;
      RECT 1.5 0.87 1.83 1.38 ;
      RECT 1.5 0.305 1.67 1.38 ;
      RECT 1.125 0.305 1.67 0.635 ;
      RECT 1.055 1.9 1.385 3.005 ;
      RECT 1.055 1.9 1.65 2.16 ;
  END
END scs130lp_a21bo_0

MACRO scs130lp_a21bo_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21bo_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.81 1.46 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.02 1.21 3.755 1.46 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 1.345 1.285 1.75 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.815 0.465 3.075 ;
        RECT 0.085 0.325 0.365 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.115 -0.085 3.445 1.04 ;
        RECT 1.725 -0.085 2.055 0.465 ;
        RECT 0.64 -0.085 0.97 0.465 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.635 1.97 2.965 3.415 ;
        RECT 0.635 2.66 0.965 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.175 1.63 3.415 3.075 ;
      RECT 2.195 1.63 2.455 3.075 ;
      RECT 2.195 1.63 3.415 1.8 ;
      RECT 1.725 2.32 2.025 3.075 ;
      RECT 1.805 1.845 2.025 3.075 ;
      RECT 0.655 2.32 2.025 2.49 ;
      RECT 0.655 0.635 0.825 2.49 ;
      RECT 0.535 1.295 0.825 1.625 ;
      RECT 2.245 0.255 2.575 1.04 ;
      RECT 0.655 0.635 2.575 0.805 ;
      RECT 1.16 1.93 1.635 2.14 ;
      RECT 1.465 0.975 1.635 2.14 ;
      RECT 1.465 1.345 1.895 1.675 ;
      RECT 1.185 0.975 1.635 1.175 ;
  END
END scs130lp_a21bo_1

MACRO scs130lp_a21bo_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21bo_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.53 1.2 3.205 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.185 3.685 1.515 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 1.21 1.455 2.12 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.61 0.325 0.825 2.155 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.415 -0.085 3.745 1.015 ;
        RECT 2.085 -0.085 2.415 0.69 ;
        RECT 0.995 -0.085 1.3 1.04 ;
        RECT 0.11 -0.085 0.44 1.205 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.965 2.025 3.295 3.415 ;
        RECT 0.97 2.665 1.3 3.415 ;
        RECT 0.11 2.665 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.465 1.685 3.745 3.075 ;
      RECT 2.53 1.685 2.795 3.075 ;
      RECT 2.53 1.685 3.745 1.855 ;
      RECT 2.085 1.815 2.36 3.075 ;
      RECT 2.185 0.86 2.36 3.075 ;
      RECT 0.11 2.325 2.36 2.495 ;
      RECT 0.11 1.375 0.44 2.495 ;
      RECT 2.185 0.86 2.845 1.03 ;
      RECT 2.585 0.255 2.845 1.03 ;
      RECT 1.625 0.795 1.885 2.155 ;
      RECT 1.625 1.055 2.015 1.625 ;
      RECT 1.625 0.795 1.915 1.625 ;
      RECT 1.495 0.795 1.915 1.04 ;
  END
END scs130lp_a21bo_2

MACRO scs130lp_a21bo_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21bo_4 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.9 1.345 5.265 1.77 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.435 1.34 6.01 1.645 ;
        RECT 4.475 1.94 5.665 2.12 ;
        RECT 5.435 1.34 5.665 2.12 ;
        RECT 4.475 1.335 4.645 2.12 ;
        RECT 4.28 1.335 4.645 1.625 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.2 0.805 1.76 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1844 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.93 2.725 2.2 ;
        RECT 0.995 1.8 2.725 2.2 ;
        RECT 0.995 1.005 2.48 1.175 ;
        RECT 2.3 0.255 2.48 1.175 ;
        RECT 1.44 0.255 1.63 1.175 ;
        RECT 0.995 1.005 1.165 2.2 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.855 -0.085 6.135 1.095 ;
        RECT 4.005 -0.085 4.335 0.825 ;
        RECT 2.67 -0.085 3.475 0.825 ;
        RECT 1.8 -0.085 2.13 0.825 ;
        RECT 0.6 -0.085 1.27 0.835 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.375 2.63 5.705 3.415 ;
        RECT 4.475 2.63 4.805 3.415 ;
        RECT 2.355 2.71 2.685 3.415 ;
        RECT 1.495 2.71 1.825 3.415 ;
        RECT 0.635 2.71 0.965 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.875 1.815 6.135 3.075 ;
      RECT 4.975 2.29 5.205 3.075 ;
      RECT 3.245 2.905 4.305 3.075 ;
      RECT 4.115 1.795 4.305 3.075 ;
      RECT 3.245 2.045 3.445 3.075 ;
      RECT 4.115 2.29 6.135 2.46 ;
      RECT 5.835 1.815 6.135 2.46 ;
      RECT 5.435 0.255 5.685 1.095 ;
      RECT 4.515 0.255 4.845 0.825 ;
      RECT 4.515 0.255 5.685 0.425 ;
      RECT 3.615 0.995 3.945 2.735 ;
      RECT 1.345 1.355 2.82 1.535 ;
      RECT 2.65 0.995 2.82 1.535 ;
      RECT 2.65 0.995 5.215 1.165 ;
      RECT 5.015 0.595 5.215 1.165 ;
      RECT 3.645 0.255 3.835 2.735 ;
      RECT 0.09 1.93 0.455 3.075 ;
      RECT 0.09 2.37 3.075 2.54 ;
      RECT 2.905 1.705 3.075 2.54 ;
      RECT 0.09 0.255 0.27 3.075 ;
      RECT 2.99 1.345 3.32 1.875 ;
      RECT 0.09 0.255 0.43 1.03 ;
  END
END scs130lp_a21bo_4

MACRO scs130lp_a21bo_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21bo_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.495 1.55 2.825 1.935 ;
        RECT 1.595 1.55 2.825 1.72 ;
        RECT 1.595 1.25 1.925 1.72 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.28 1.355 1.78 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.035 3.335 1.78 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 2.025 0.495 3.065 ;
        RECT 0.09 0.265 0.445 0.715 ;
        RECT 0.09 0.265 0.26 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.515 -0.085 2.845 0.505 ;
        RECT 0.905 -0.085 1.235 0.715 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.855 2.115 3.185 3.415 ;
        RECT 0.695 2.31 1.025 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.385 2.075 3.715 3.065 ;
      RECT 3.545 0.685 3.715 3.065 ;
      RECT 2.25 0.685 2.58 1.135 ;
      RECT 2.25 0.685 3.715 0.855 ;
      RECT 3.305 0.265 3.635 0.855 ;
      RECT 1.235 2.895 2.655 3.065 ;
      RECT 2.325 2.115 2.655 3.065 ;
      RECT 1.235 2.31 1.565 3.065 ;
      RECT 1.765 1.96 2.095 2.715 ;
      RECT 0.675 1.96 2.095 2.13 ;
      RECT 0.675 0.895 0.845 2.13 ;
      RECT 0.44 0.895 0.845 1.565 ;
      RECT 0.44 0.895 2.055 1.065 ;
      RECT 1.725 0.265 2.055 1.065 ;
  END
END scs130lp_a21bo_lp

MACRO scs130lp_a21bo_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21bo_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.765 2.445 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.975 0.84 3.205 1.75 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.025 1.285 2.12 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.685 0.365 3.015 ;
        RECT 0.155 0.47 0.365 0.8 ;
        RECT 0.155 0.47 0.325 3.015 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.975 -0.085 3.165 0.545 ;
        RECT 1.53 -0.085 1.86 0.485 ;
        RECT 0.585 -0.085 0.795 0.8 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.56 2.325 2.77 3.415 ;
        RECT 0.585 2.755 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.99 1.975 3.2 2.505 ;
      RECT 2.13 1.975 2.34 2.505 ;
      RECT 2.13 1.975 3.2 2.145 ;
      RECT 0.505 2.335 1.91 2.505 ;
      RECT 1.7 1.625 1.91 2.505 ;
      RECT 0.505 1.475 0.675 2.505 ;
      RECT 1.7 1.625 2.795 1.795 ;
      RECT 2.625 0.285 2.795 1.795 ;
      RECT 2.04 0.285 2.795 0.495 ;
      RECT 1.705 0.675 1.875 1.435 ;
      RECT 1.015 0.675 1.875 0.845 ;
      RECT 1.015 0.515 1.225 0.845 ;
      RECT 1.015 2.695 1.735 3.025 ;
  END
END scs130lp_a21bo_m

MACRO scs130lp_a21boi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21boi_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.72 0.78 2.255 1.875 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 0.78 2.795 1.855 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 1.565 0.9 2.5 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2872 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.315 0.28 1.625 0.61 ;
        RECT 1.07 1.565 1.485 3.065 ;
        RECT 1.315 0.28 1.485 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.085 -0.085 2.415 0.61 ;
        RECT 0.55 -0.085 1.145 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.055 2.405 2.32 3.415 ;
        RECT 0.525 2.67 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.49 2.055 2.785 3.065 ;
      RECT 1.655 2.055 1.885 3.065 ;
      RECT 1.655 2.055 2.785 2.225 ;
      RECT 0.095 0.28 0.355 3 ;
      RECT 0.095 0.78 1.09 1.395 ;
      RECT 0.095 0.28 0.38 1.395 ;
  END
END scs130lp_a21boi_0

MACRO scs130lp_a21boi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21boi_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.83 0.375 2.275 1.015 ;
        RECT 1.83 0.375 2.255 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.185 2.795 1.515 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.785 0.355 2.13 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6237 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.095 1.21 1.66 1.515 ;
        RECT 1.415 0.255 1.66 1.515 ;
        RECT 1.095 1.21 1.355 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.445 -0.085 2.775 1.015 ;
        RECT 1 -0.085 1.245 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.97 2.025 2.3 3.415 ;
        RECT 0.525 2.64 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.47 1.685 2.775 3.075 ;
      RECT 1.525 1.685 1.8 3.075 ;
      RECT 1.525 1.685 2.775 1.855 ;
      RECT 0.095 2.3 0.355 2.915 ;
      RECT 0.095 2.3 0.925 2.47 ;
      RECT 0.66 1.345 0.925 2.47 ;
      RECT 0.66 0.28 0.83 2.47 ;
      RECT 0.425 0.28 0.83 0.61 ;
  END
END scs130lp_a21boi_1

MACRO scs130lp_a21boi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21boi_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.79 1.425 3.315 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.515 1.355 4.06 1.645 ;
        RECT 2.425 1.925 3.745 2.12 ;
        RECT 3.515 1.355 3.745 2.12 ;
        RECT 2.425 1.425 2.595 2.12 ;
        RECT 2.25 1.425 2.595 1.595 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.32 0.47 2.49 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8904 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.075 3.325 1.245 ;
        RECT 2.995 0.605 3.325 1.245 ;
        RECT 1.545 1.82 1.875 2.73 ;
        RECT 1.545 0.285 1.805 1.245 ;
        RECT 1.545 0.285 1.795 2.73 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.89 -0.085 4.185 1.185 ;
        RECT 1.975 -0.085 2.305 0.905 ;
        RECT 1.115 -0.085 1.375 1.17 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.425 2.63 3.755 3.415 ;
        RECT 2.485 2.64 2.815 3.415 ;
        RECT 0.14 2.66 0.47 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.925 1.815 4.185 3.075 ;
      RECT 1.115 2.905 2.315 3.075 ;
      RECT 2.045 2.29 2.315 3.075 ;
      RECT 2.985 2.29 3.255 2.97 ;
      RECT 1.115 1.83 1.375 3.075 ;
      RECT 2.045 2.29 4.185 2.46 ;
      RECT 3.915 1.815 4.185 2.46 ;
      RECT 2.045 1.83 2.245 3.075 ;
      RECT 3.495 0.265 3.72 1.185 ;
      RECT 2.485 0.265 2.815 0.905 ;
      RECT 2.485 0.265 3.72 0.435 ;
      RECT 0.64 0.37 0.9 2.875 ;
      RECT 0.64 1.34 1.165 1.605 ;
      RECT 0.64 0.37 0.92 1.605 ;
  END
END scs130lp_a21boi_2

MACRO scs130lp_a21boi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21boi_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 1.415 5.165 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.335 1.21 6.605 1.515 ;
        RECT 3.03 1.075 5.605 1.245 ;
        RECT 3.03 1.075 3.315 1.515 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.805 1.75 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.135 0.695 4.885 0.895 ;
        RECT 2.545 0.695 2.86 1.75 ;
        RECT 2.435 1.715 2.725 2.665 ;
        RECT 1.315 1.035 2.86 1.205 ;
        RECT 2.135 0.695 2.86 1.205 ;
        RECT 1.505 1.715 2.725 2.035 ;
        RECT 2.135 0.255 2.365 1.205 ;
        RECT 1.505 1.715 1.765 2.485 ;
        RECT 1.315 0.37 1.485 1.205 ;
        RECT 1.275 0.37 1.485 0.7 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 6.305 -0.085 6.605 1.04 ;
        RECT 5.485 -0.085 5.715 0.565 ;
        RECT 2.535 -0.085 3.095 0.525 ;
        RECT 1.655 -0.085 1.965 0.865 ;
        RECT 0.775 -0.085 1.105 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.845 2.105 6.175 3.415 ;
        RECT 4.985 2.26 5.315 3.415 ;
        RECT 3.265 2.26 4.455 2.495 ;
        RECT 3.265 2.26 3.595 3.415 ;
        RECT 0.555 2.26 0.885 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.345 1.685 6.605 3.075 ;
      RECT 5.485 1.685 5.665 3.075 ;
      RECT 1.075 2.835 3.095 3.075 ;
      RECT 2.895 1.92 3.095 3.075 ;
      RECT 3.765 2.665 4.815 3.065 ;
      RECT 4.625 1.92 4.815 3.065 ;
      RECT 1.075 2.665 2.265 3.075 ;
      RECT 1.935 2.205 2.265 3.075 ;
      RECT 1.075 2.26 1.335 3.075 ;
      RECT 2.895 1.92 5.665 2.09 ;
      RECT 5.335 1.685 6.605 1.925 ;
      RECT 5.905 0.255 6.135 1.04 ;
      RECT 5.055 0.735 6.135 0.905 ;
      RECT 5.885 0.255 6.135 0.905 ;
      RECT 5.055 0.255 5.315 0.905 ;
      RECT 3.265 0.255 5.315 0.525 ;
      RECT 0.125 1.92 0.385 3.075 ;
      RECT 0.125 1.92 1.195 2.09 ;
      RECT 0.975 1.375 1.195 2.09 ;
      RECT 0.975 1.375 2.375 1.545 ;
      RECT 0.975 0.87 1.145 2.09 ;
      RECT 0.325 0.87 1.145 1.04 ;
      RECT 0.325 0.255 0.605 1.04 ;
  END
END scs130lp_a21boi_4

MACRO scs130lp_a21boi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21boi_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.46 1.315 1.79 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.81 0.835 1.14 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.825 2.855 1.495 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.695 2.025 2.045 3.065 ;
        RECT 1.495 1.92 1.865 2.15 ;
        RECT 1.495 0.265 1.665 2.15 ;
        RECT 1.225 0.265 1.665 0.675 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.015 -0.085 2.345 0.675 ;
        RECT 0.405 -0.085 0.735 0.63 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.37 2.025 2.7 3.415 ;
        RECT 0.655 2.68 0.985 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.9 1.675 3.23 3.065 ;
      RECT 3.06 0.265 3.23 3.065 ;
      RECT 2.045 1.675 3.23 1.845 ;
      RECT 1.845 1.07 2.215 1.74 ;
      RECT 2.9 0.265 3.23 0.645 ;
      RECT 1.185 2.33 1.515 3.065 ;
      RECT 0.125 2.025 0.455 3.065 ;
      RECT 0.125 2.33 1.515 2.5 ;
  END
END scs130lp_a21boi_lp

MACRO scs130lp_a21boi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21boi_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 0.47 1.765 1.475 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.765 2.38 1.435 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.48 0.805 0.805 2.12 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.265 1.345 2.285 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.11 -0.085 2.44 0.485 ;
        RECT 0.725 -0.085 0.935 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.935 2.145 2.265 3.415 ;
        RECT 0.525 2.845 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.445 1.795 2.635 2.285 ;
      RECT 1.565 1.795 1.755 2.285 ;
      RECT 1.565 1.795 2.635 1.965 ;
      RECT 1.055 2.495 1.225 3.065 ;
      RECT 0.13 2.495 0.345 2.985 ;
      RECT 0.13 2.495 1.225 2.665 ;
      RECT 0.13 0.295 0.3 2.985 ;
      RECT 0.13 0.295 0.505 0.625 ;
  END
END scs130lp_a21boi_m

MACRO scs130lp_a21o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21o_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.955 0.78 2.31 1.835 ;
        RECT 1.955 0.38 2.3 1.835 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.48 0.78 2.795 1.83 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.385 1.08 1.785 1.83 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.28 0.88 0.61 ;
        RECT 0.085 0.28 0.395 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.47 -0.085 2.72 0.61 ;
        RECT 1.05 -0.085 1.38 0.57 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.04 2.345 2.295 3.415 ;
        RECT 0.565 2.395 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.465 2.005 2.76 3.025 ;
      RECT 1.595 2.005 1.87 3.025 ;
      RECT 1.595 2.005 2.76 2.175 ;
      RECT 1.14 2.055 1.425 3.025 ;
      RECT 1.035 0.74 1.205 2.225 ;
      RECT 0.71 0.78 1.205 1.525 ;
      RECT 1.55 0.28 1.785 0.91 ;
      RECT 1.035 0.74 1.785 0.91 ;
  END
END scs130lp_a21o_0

MACRO scs130lp_a21o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21o_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.74 1.185 2.255 1.515 ;
        RECT 1.94 0.34 2.255 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.185 2.795 1.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.345 1.385 1.75 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 0.255 0.355 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.435 -0.085 2.765 1.015 ;
        RECT 0.53 -0.085 1.22 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.96 2.025 2.29 3.415 ;
        RECT 0.525 2.27 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.46 1.685 2.765 3.075 ;
      RECT 1.555 1.685 1.745 3.075 ;
      RECT 1.555 1.685 2.765 1.855 ;
      RECT 1.045 1.92 1.315 3.075 ;
      RECT 0.715 1.92 1.315 2.1 ;
      RECT 0.715 0.985 0.885 2.1 ;
      RECT 0.525 1.185 0.885 1.515 ;
      RECT 0.715 0.985 1.57 1.155 ;
      RECT 1.39 0.255 1.72 1.015 ;
  END
END scs130lp_a21o_1

MACRO scs130lp_a21o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21o_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 0.315 2.735 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.185 3.27 1.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.345 1.82 1.76 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.795 0.255 0.985 1.155 ;
        RECT 0.585 0.985 0.815 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.905 -0.085 3.175 1.015 ;
        RECT 1.155 -0.085 1.485 0.815 ;
        RECT 0.295 -0.085 0.625 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.385 2.025 2.715 3.415 ;
        RECT 0.985 2.27 1.315 3.415 ;
        RECT 0.125 1.815 0.415 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.885 1.685 3.105 3.075 ;
      RECT 1.99 1.685 2.215 3.075 ;
      RECT 1.99 1.685 3.105 1.855 ;
      RECT 1.505 1.93 1.82 3.075 ;
      RECT 0.985 1.93 1.82 2.1 ;
      RECT 0.985 1.345 1.325 2.1 ;
      RECT 1.155 0.985 1.325 2.1 ;
      RECT 1.155 0.985 1.895 1.155 ;
      RECT 1.705 0.255 1.895 1.155 ;
  END
END scs130lp_a21o_2

MACRO scs130lp_a21o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21o_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.265 1.21 4.645 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.955 1.345 5.43 1.645 ;
        RECT 3.915 1.95 5.125 2.12 ;
        RECT 4.955 1.345 5.125 2.12 ;
        RECT 3.915 1.295 4.085 2.12 ;
        RECT 3.7 1.295 4.085 1.625 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 2.935 1.76 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.075 2.035 1.245 ;
        RECT 1.845 0.255 2.035 1.245 ;
        RECT 1.725 1.78 1.915 3.075 ;
        RECT 0.155 1.78 1.915 1.985 ;
        RECT 0.985 0.255 1.175 1.245 ;
        RECT 0.865 1.78 1.055 3.075 ;
        RECT 0.155 1.075 0.805 1.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 5.26 -0.085 5.555 1.105 ;
        RECT 3.475 -0.085 3.815 0.69 ;
        RECT 2.24 -0.085 2.895 0.7 ;
        RECT 1.345 -0.085 1.675 0.905 ;
        RECT 0.485 -0.085 0.815 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.795 2.64 5.125 3.415 ;
        RECT 3.915 2.64 4.245 3.415 ;
        RECT 2.085 1.815 2.385 3.415 ;
        RECT 1.225 2.155 1.555 3.415 ;
        RECT 0.365 2.155 0.695 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.295 1.815 5.495 3.075 ;
      RECT 4.415 2.3 4.625 3.075 ;
      RECT 2.605 2.905 3.735 3.075 ;
      RECT 3.535 1.815 3.735 3.075 ;
      RECT 2.605 1.93 2.865 3.075 ;
      RECT 3.535 2.3 5.495 2.47 ;
      RECT 3.535 1.815 3.745 2.47 ;
      RECT 4.795 0.255 5.09 1.105 ;
      RECT 3.985 0.255 4.235 0.69 ;
      RECT 3.985 0.255 5.09 0.435 ;
      RECT 3.035 1.91 3.365 2.735 ;
      RECT 3.105 0.86 3.365 2.735 ;
      RECT 0.985 1.415 2.375 1.61 ;
      RECT 2.205 0.87 2.375 1.61 ;
      RECT 2.205 0.87 3.365 1.04 ;
      RECT 3.065 0.255 3.305 1.04 ;
      RECT 4.405 0.605 4.625 1.03 ;
      RECT 3.065 0.86 4.625 1.03 ;
  END
END scs130lp_a21o_4

MACRO scs130lp_a21o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21o_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.94 1.125 1.315 1.795 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.55 1.78 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.51 1.125 1.84 1.795 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.915 0.265 3.245 3 ;
        RECT 2.815 0.265 3.245 1.78 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.995 -0.085 2.325 0.595 ;
        RECT 0.245 -0.085 0.575 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.385 1.96 2.715 3.415 ;
        RECT 0.675 2.325 1.005 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.735 2.025 2.19 3.065 ;
      RECT 2.02 0.775 2.19 3.065 ;
      RECT 2.02 0.775 2.63 1.485 ;
      RECT 1.205 0.775 2.63 0.945 ;
      RECT 1.205 0.265 1.535 0.945 ;
      RECT 1.205 1.975 1.535 3.065 ;
      RECT 0.145 1.975 0.475 3.065 ;
      RECT 0.145 1.975 1.535 2.145 ;
  END
END scs130lp_a21o_lp

MACRO scs130lp_a21o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21o_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.8 0.84 2.245 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.47 2.725 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.07 1.21 1.285 2.12 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.345 0.635 0.675 ;
        RECT 0.155 0.345 0.345 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.015 -0.085 2.345 0.485 ;
        RECT 0.855 -0.085 1.065 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.085 2.65 2.295 3.415 ;
        RECT 0.525 2.845 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.515 2.3 2.725 2.85 ;
      RECT 1.655 2.3 1.865 2.85 ;
      RECT 1.655 2.3 2.725 2.47 ;
      RECT 1.225 2.345 1.435 2.85 ;
      RECT 0.525 2.345 1.435 2.515 ;
      RECT 0.525 0.86 0.695 2.515 ;
      RECT 0.525 0.86 1.495 1.03 ;
      RECT 1.285 0.33 1.495 1.03 ;
  END
END scs130lp_a21o_m

MACRO scs130lp_a21oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21oi_0 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 0.74 0.925 1.835 ;
        RECT 0.625 0.395 0.925 1.835 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.4 1.835 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.455 0.78 1.83 1.395 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2872 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.51 1.565 1.835 3.025 ;
        RECT 1.095 1.565 1.835 1.75 ;
        RECT 1.095 0.28 1.34 0.61 ;
        RECT 1.095 0.28 1.285 1.75 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.51 -0.085 1.805 0.61 ;
        RECT 0.205 -0.085 0.455 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.645 2.345 0.915 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.085 2.005 1.34 3.025 ;
      RECT 0.185 2.005 0.475 3.025 ;
      RECT 0.185 2.005 1.34 2.175 ;
  END
END scs130lp_a21oi_0

MACRO scs130lp_a21oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21oi_1 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.345 1.02 1.75 ;
        RECT 0.625 0.37 0.815 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.455 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.21 1.835 1.78 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6615 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.95 1.835 3.075 ;
        RECT 1.19 1.95 1.835 2.13 ;
        RECT 1.19 0.325 1.36 2.13 ;
        RECT 0.985 0.325 1.36 1.165 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.53 -0.085 1.81 1.04 ;
        RECT 0.095 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.56 2.64 0.89 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.06 2.3 1.355 3.075 ;
      RECT 0.095 1.93 0.39 3.075 ;
      RECT 0.095 2.3 1.355 2.47 ;
      RECT 0.095 1.93 1.02 2.47 ;
  END
END scs130lp_a21oi_1

MACRO scs130lp_a21oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21oi_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.205 1.355 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.345 1.87 1.675 ;
        RECT 0.125 1.605 1.765 1.785 ;
        RECT 0.125 1.295 0.455 1.785 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.04 1.425 2.8 1.76 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8232 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.285 1.93 3.275 2.1 ;
        RECT 2.97 1.005 3.275 2.1 ;
        RECT 2.345 1.005 3.275 1.175 ;
        RECT 2.285 1.93 2.615 2.735 ;
        RECT 1.025 0.865 2.545 1.035 ;
        RECT 2.335 0.255 2.545 1.035 ;
        RECT 1.025 0.595 1.26 1.035 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.715 -0.085 3.045 0.835 ;
        RECT 1.835 -0.085 2.165 0.695 ;
        RECT 0.095 -0.085 0.355 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.405 2.295 1.735 3.415 ;
        RECT 0.525 2.295 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.905 2.905 3.045 3.075 ;
      RECT 2.785 2.27 3.045 3.075 ;
      RECT 1.025 1.955 1.235 3.075 ;
      RECT 0.095 1.955 0.355 3.075 ;
      RECT 1.905 1.955 2.115 3.075 ;
      RECT 0.095 1.955 2.115 2.125 ;
      RECT 0.525 0.255 0.855 1.035 ;
      RECT 1.43 0.255 1.665 0.695 ;
      RECT 0.525 0.255 1.665 0.425 ;
  END
END scs130lp_a21oi_2

MACRO scs130lp_a21oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21oi_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.2 3.23 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.615 3.675 1.785 ;
        RECT 3.4 1.345 3.675 1.785 ;
        RECT 0.105 1.375 1.765 1.785 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.885 1.425 5.235 1.76 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.055 1.93 5.585 2.1 ;
        RECT 5.415 1.085 5.585 2.1 ;
        RECT 4.07 1.085 5.585 1.255 ;
        RECT 4.91 1.93 5.155 2.735 ;
        RECT 4.94 0.255 5.13 1.255 ;
        RECT 4.055 1.93 4.295 2.735 ;
        RECT 4.07 0.255 4.26 1.255 ;
        RECT 1.82 0.82 4.26 1.03 ;
        RECT 4.06 0.255 4.26 1.03 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 5.3 -0.085 5.63 0.915 ;
        RECT 4.44 -0.085 4.77 0.915 ;
        RECT 3.56 -0.085 3.89 0.65 ;
        RECT 0.96 -0.085 1.29 0.865 ;
        RECT 0.1 -0.085 0.39 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 3.11 2.295 3.44 3.415 ;
        RECT 2.25 2.295 2.58 3.415 ;
        RECT 1.39 2.295 1.72 3.415 ;
        RECT 0.53 2.295 0.86 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.61 2.905 5.63 3.075 ;
      RECT 5.325 2.27 5.63 3.075 ;
      RECT 2.75 1.955 2.94 3.075 ;
      RECT 1.9 1.955 2.08 3.075 ;
      RECT 1.03 1.955 1.22 3.075 ;
      RECT 0.1 1.955 0.36 3.075 ;
      RECT 4.465 2.27 4.74 3.075 ;
      RECT 3.61 1.955 3.885 3.075 ;
      RECT 0.1 1.955 3.885 2.125 ;
      RECT 0.56 1.035 1.65 1.205 ;
      RECT 1.46 0.255 1.65 1.205 ;
      RECT 0.56 0.255 0.79 1.205 ;
      RECT 1.46 0.255 3.38 0.64 ;
  END
END scs130lp_a21oi_4

MACRO scs130lp_a21oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21oi_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.9 1.075 1.315 1.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.855 0.55 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.075 1.825 1.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4614 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.725 2.025 2.275 3.065 ;
        RECT 2.075 0.725 2.275 3.065 ;
        RECT 1.165 0.725 2.275 0.895 ;
        RECT 1.165 0.265 1.495 0.895 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.955 -0.085 2.285 0.545 ;
        RECT 0.205 -0.085 0.535 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.665 2.275 0.995 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.195 1.925 1.525 3.065 ;
      RECT 0.135 1.925 0.465 3.065 ;
      RECT 0.135 1.925 1.525 2.095 ;
  END
END scs130lp_a21oi_lp

MACRO scs130lp_a21oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a21oi_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 0.9 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.36 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.08 1.47 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2604 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.445 2.53 1.82 2.86 ;
        RECT 1.65 0.665 1.82 2.86 ;
        RECT 1.08 0.665 1.82 0.835 ;
        RECT 1.08 0.345 1.25 0.835 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.43 -0.085 1.76 0.485 ;
        RECT 0.195 -0.085 0.405 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.585 2.65 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.155 2.3 0.365 2.83 ;
      RECT 1.015 2.3 1.225 2.81 ;
      RECT 0.155 2.3 1.225 2.47 ;
  END
END scs130lp_a21oi_m

MACRO scs130lp_a221o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221o_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.54 0.84 1.845 1.605 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.9 1.065 1.36 1.615 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 0.84 2.27 1.51 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.495 1.05 2.84 1.585 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.36 0.995 3.755 1.665 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 0.28 0.535 0.555 ;
        RECT 0.09 2.4 0.475 3.075 ;
        RECT 0.09 0.28 0.335 1.39 ;
        RECT 0.09 0.28 0.27 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.78 -0.085 3.11 0.475 ;
        RECT 0.715 -0.085 1.03 0.555 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.52 2.4 1.815 3.415 ;
        RECT 0.645 2.4 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.455 1.845 3.715 2.795 ;
      RECT 0.44 1.56 0.675 2.23 ;
      RECT 0.505 0.725 0.675 2.23 ;
      RECT 3.01 1.845 3.715 2.015 ;
      RECT 3.01 0.645 3.19 2.015 ;
      RECT 0.505 0.725 1.37 0.895 ;
      RECT 1.2 0.28 1.37 0.895 ;
      RECT 2.44 0.645 3.575 0.815 ;
      RECT 3.28 0.28 3.575 0.815 ;
      RECT 2.44 0.28 2.61 0.815 ;
      RECT 1.2 0.28 2.61 0.61 ;
      RECT 2.005 2.905 3.285 3.075 ;
      RECT 2.955 2.185 3.285 3.075 ;
      RECT 2.005 2.135 2.285 3.075 ;
      RECT 1.095 1.785 1.35 3.075 ;
      RECT 2.455 1.785 2.785 2.735 ;
      RECT 1.095 1.785 2.785 1.955 ;
  END
END scs130lp_a221o_0

MACRO scs130lp_a221o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221o_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.185 1.855 1.515 ;
        RECT 1.535 0.33 1.765 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.185 1.365 1.515 ;
        RECT 1.115 0.33 1.365 1.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.385 1.185 2.785 1.515 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.955 1.185 3.29 1.515 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.46 1.185 4.235 1.435 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.255 0.425 1.075 ;
        RECT 0.085 0.255 0.345 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.13 -0.085 3.46 0.665 ;
        RECT 0.615 -0.085 0.945 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 1.73 2.365 2.06 3.415 ;
        RECT 0.525 2.025 1.195 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.64 1.685 3.97 3.075 ;
      RECT 0.515 1.685 3.97 1.855 ;
      RECT 2.025 0.255 2.205 1.855 ;
      RECT 0.515 1.305 0.765 1.855 ;
      RECT 1.935 0.835 3.97 1.015 ;
      RECT 3.7 0.255 3.97 1.015 ;
      RECT 1.935 0.255 2.58 1.015 ;
      RECT 2.25 2.905 3.47 3.075 ;
      RECT 3.25 2.025 3.47 3.075 ;
      RECT 2.25 2.365 2.58 3.075 ;
      RECT 1.365 2.025 1.56 3.075 ;
      RECT 2.75 2.025 3.08 2.735 ;
      RECT 1.365 2.025 3.08 2.195 ;
  END
END scs130lp_a221o_1

MACRO scs130lp_a221o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221o_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.425 2.405 2.26 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.445 1.425 1.835 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 1.425 3.805 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.995 1.21 4.645 1.75 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 1.425 3.265 1.76 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 0.255 0.815 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.14 -0.085 4.47 1.04 ;
        RECT 2.81 -0.085 3.14 0.905 ;
        RECT 0.985 -0.085 1.655 0.905 ;
        RECT 0.125 -0.085 0.425 1.125 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 2.11 2.845 2.44 3.415 ;
        RECT 1.105 1.92 1.435 3.415 ;
        RECT 0.125 1.815 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.24 2.77 4.47 3.075 ;
      RECT 4.17 1.92 4.47 3.075 ;
      RECT 1.645 2.43 1.94 3.075 ;
      RECT 1.645 2.43 4 2.6 ;
      RECT 3.67 1.92 4 2.6 ;
      RECT 1.645 1.92 1.905 3.075 ;
      RECT 2.585 1.93 3.08 2.26 ;
      RECT 2.585 1.075 2.755 2.26 ;
      RECT 0.985 1.075 1.235 1.545 ;
      RECT 2.585 1.075 3.57 1.255 ;
      RECT 3.31 0.255 3.57 1.255 ;
      RECT 0.985 1.075 3.57 1.245 ;
      RECT 2.115 0.255 2.445 1.245 ;
  END
END scs130lp_a221o_2

MACRO scs130lp_a221o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221o_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.375 1.185 3.955 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.19 1.185 3.205 1.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.295 1.195 6.135 1.525 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.64 1.405 7.525 1.75 ;
        RECT 6.63 1.405 7.525 1.62 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.465 1.195 5.125 1.525 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.47 1.755 1.66 3.075 ;
        RECT 0.11 1.06 1.66 1.23 ;
        RECT 1.47 0.255 1.66 1.23 ;
        RECT 0.11 1.755 1.66 1.925 ;
        RECT 0.61 1.045 1.66 1.23 ;
        RECT 0.61 0.255 0.8 1.23 ;
        RECT 0.61 1.755 0.79 3.075 ;
        RECT 0.11 1.06 0.335 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.74 -0.085 7.07 0.895 ;
        RECT 4.535 -0.085 4.795 0.685 ;
        RECT 2.69 -0.085 3.02 0.675 ;
        RECT 1.83 -0.085 2.16 1.015 ;
        RECT 0.97 -0.085 1.3 0.875 ;
        RECT 0.11 -0.085 0.44 0.89 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 3.55 2.385 3.88 3.415 ;
        RECT 2.69 2.395 3.02 3.415 ;
        RECT 1.83 2.045 2.16 3.415 ;
        RECT 0.97 2.095 1.3 3.415 ;
        RECT 0.11 2.095 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.37 1.065 7.5 1.235 ;
      RECT 7.24 0.255 7.5 1.235 ;
      RECT 6.37 0.255 6.57 1.235 ;
      RECT 5.405 0.685 6.57 1.015 ;
      RECT 6.31 0.255 6.57 1.015 ;
      RECT 4.07 2.895 6.98 3.065 ;
      RECT 6.65 1.92 6.98 3.065 ;
      RECT 4.07 2.785 6.12 3.065 ;
      RECT 5.79 2.055 6.12 3.065 ;
      RECT 2.33 2.045 2.52 3.075 ;
      RECT 3.19 2.045 3.38 3.065 ;
      RECT 6.29 1.705 6.47 2.725 ;
      RECT 4.07 2.445 5.62 2.615 ;
      RECT 5.36 1.705 5.62 2.615 ;
      RECT 4.07 2.045 4.315 2.615 ;
      RECT 2.33 2.045 3.38 2.225 ;
      RECT 2.33 2.045 4.315 2.215 ;
      RECT 5.36 1.705 6.47 1.875 ;
      RECT 4.5 1.705 4.83 2.275 ;
      RECT 1.85 1.705 4.83 1.875 ;
      RECT 1.85 1.69 4.295 1.875 ;
      RECT 4.125 0.255 4.295 1.875 ;
      RECT 1.85 1.4 2.02 1.875 ;
      RECT 0.505 1.4 2.02 1.585 ;
      RECT 4.125 0.855 5.235 1.025 ;
      RECT 4.965 0.255 5.235 1.025 ;
      RECT 4.125 0.255 4.365 1.025 ;
      RECT 3.21 0.255 3.53 0.675 ;
      RECT 4.965 0.255 6.12 0.515 ;
      RECT 3.21 0.255 4.365 0.425 ;
      RECT 2.33 0.845 3.955 1.015 ;
      RECT 3.7 0.595 3.955 1.015 ;
      RECT 2.33 0.255 2.52 1.015 ;
  END
END scs130lp_a221o_4

MACRO scs130lp_a221o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221o_lp 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.93 0.44 2.275 1.53 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.07 1.265 1.4 1.935 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.5 1.18 2.83 1.51 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.18 3.715 1.78 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 1.17 4.36 1.84 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.92 0.835 3.065 ;
        RECT 0.125 0.565 0.685 0.735 ;
        RECT 0.355 0.31 0.685 0.735 ;
        RECT 0.125 0.565 0.295 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.275 -0.085 3.605 0.64 ;
        RECT 1.225 -0.085 1.555 0.735 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 2.115 2.41 2.445 3.415 ;
        RECT 1.015 2.115 1.345 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.295 2.02 4.71 3.02 ;
      RECT 4.54 0.31 4.71 3.02 ;
      RECT 1.58 1.71 3.18 1.88 ;
      RECT 3.01 0.82 3.18 1.88 ;
      RECT 1.58 0.915 1.75 1.88 ;
      RECT 0.48 0.915 0.81 1.585 ;
      RECT 0.48 0.915 1.75 1.085 ;
      RECT 2.455 0.82 4.71 0.99 ;
      RECT 4.155 0.31 4.71 0.99 ;
      RECT 2.455 0.31 2.785 0.99 ;
      RECT 2.705 2.895 4.095 3.065 ;
      RECT 3.765 2.02 4.095 3.065 ;
      RECT 2.705 2.41 3.035 3.065 ;
      RECT 1.585 2.06 1.915 3.065 ;
      RECT 3.235 2.06 3.565 2.715 ;
      RECT 1.585 2.06 3.565 2.23 ;
  END
END scs130lp_a221o_lp

MACRO scs130lp_a221o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221o_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.47 1.44 1.095 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 0.805 1.485 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.97 1.155 2.245 1.485 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.43 1.21 2.76 1.405 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 2.69 3.205 3.075 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.655 0.55 2.985 ;
        RECT 0.155 0.345 0.345 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.33 -0.085 2.66 0.485 ;
        RECT 0.525 -0.085 0.855 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.57 2.845 1.9 3.415 ;
        RECT 0.77 2.785 0.98 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.525 1.695 0.695 2.365 ;
      RECT 2.995 0.405 3.245 2.295 ;
      RECT 0.525 1.695 1.155 1.865 ;
      RECT 0.985 1.395 1.155 1.865 ;
      RECT 0.985 1.395 1.79 1.565 ;
      RECT 1.62 0.345 1.79 1.565 ;
      RECT 1.62 0.665 3.245 0.835 ;
      RECT 2.915 0.405 3.245 0.835 ;
      RECT 1.62 0.345 1.81 0.835 ;
      RECT 2.565 1.745 2.775 2.295 ;
      RECT 1.705 1.745 1.915 2.295 ;
      RECT 1.705 1.745 2.775 1.915 ;
      RECT 1.2 2.495 1.39 2.985 ;
      RECT 1.2 2.495 2.345 2.665 ;
      RECT 2.135 2.095 2.345 2.665 ;
  END
END scs130lp_a221o_m

MACRO scs130lp_a221oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221oi_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.185 1.895 1.965 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.185 2.58 1.965 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.75 0.78 3.205 1.965 ;
        RECT 1.35 0.78 3.205 1.015 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.99 1.185 1.375 1.965 ;
        RECT 0.99 1.18 1.305 1.965 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.53 1.18 0.82 2.05 ;
        RECT 0.53 1.18 0.805 2.12 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4321 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 0.28 1.905 0.61 ;
        RECT 0.155 0.78 1.17 1.01 ;
        RECT 1 0.28 1.17 1.01 ;
        RECT 0.155 2.415 0.655 3.075 ;
        RECT 0.155 0.28 0.39 1.01 ;
        RECT 0.155 0.28 0.36 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.405 -0.085 2.735 0.61 ;
        RECT 0.61 -0.085 0.83 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.815 2.825 2.145 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.815 2.135 3.145 3.075 ;
      RECT 0.825 2.305 1.145 3.075 ;
      RECT 0.975 2.135 3.145 2.305 ;
      RECT 2.315 2.475 2.645 3.075 ;
      RECT 1.315 2.475 1.645 3.075 ;
      RECT 1.315 2.475 2.645 2.655 ;
  END
END scs130lp_a221oi_0

MACRO scs130lp_a221oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221oi_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.31 1.185 2.735 1.515 ;
        RECT 2.45 0.325 2.735 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.185 3.275 1.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.21 2.04 1.515 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 1.185 1.39 1.515 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 1.21 0.86 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8841 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 0.845 2.22 1.015 ;
        RECT 1.89 0.255 2.22 1.015 ;
        RECT 0.09 0.265 0.52 1.015 ;
        RECT 0.09 0.265 0.375 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.915 -0.085 3.245 1.015 ;
        RECT 0.69 -0.085 1.375 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.44 2.045 2.77 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.975 1.705 3.245 3.075 ;
      RECT 1.95 1.705 2.27 3.075 ;
      RECT 1.045 1.705 1.375 2.735 ;
      RECT 1.045 1.705 3.245 1.875 ;
      RECT 0.545 2.905 1.78 3.075 ;
      RECT 1.545 2.045 1.78 3.075 ;
      RECT 0.545 1.92 0.855 3.075 ;
  END
END scs130lp_a221oi_1

MACRO scs130lp_a221oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221oi_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.96 1.21 5.165 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.54 1.615 5.675 1.785 ;
        RECT 5.335 1.21 5.675 1.785 ;
        RECT 3.54 1.345 3.79 1.785 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.21 2.815 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.615 3.33 1.785 ;
        RECT 3 1.375 3.33 1.785 ;
        RECT 1.025 1.425 2.255 1.785 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.465 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0584 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.785 4.465 1.04 ;
        RECT 4.205 0.665 4.465 1.04 ;
        RECT 0.635 0.255 0.895 1.04 ;
        RECT 0.525 1.92 0.855 2.735 ;
        RECT 0.635 0.255 0.855 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 5.135 -0.085 5.395 1.04 ;
        RECT 3.26 -0.085 3.59 0.615 ;
        RECT 1.065 -0.085 1.775 0.615 ;
        RECT 0.205 -0.085 0.465 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.635 2.295 4.965 3.415 ;
        RECT 3.72 2.295 4.05 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.145 1.955 5.395 3.075 ;
      RECT 4.22 1.955 4.455 3.075 ;
      RECT 1.475 2.905 3.55 3.075 ;
      RECT 3.265 1.955 3.55 3.075 ;
      RECT 2.405 2.295 2.595 3.075 ;
      RECT 1.475 2.295 1.735 3.075 ;
      RECT 3.265 1.955 5.395 2.125 ;
      RECT 4.635 0.255 4.965 1.04 ;
      RECT 3.775 0.255 4.965 0.485 ;
      RECT 0.095 2.905 1.285 3.075 ;
      RECT 1.025 1.955 1.285 3.075 ;
      RECT 0.095 1.925 0.355 3.075 ;
      RECT 2.765 1.955 3.095 2.735 ;
      RECT 1.905 1.955 2.235 2.735 ;
      RECT 1.025 1.955 3.095 2.125 ;
      RECT 1.955 0.285 3.085 0.615 ;
  END
END scs130lp_a221oi_2

MACRO scs130lp_a221oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221oi_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.83 1.2 8.075 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.245 1.21 9.995 1.435 ;
        RECT 6.41 1.615 8.485 1.785 ;
        RECT 8.245 1.21 8.485 1.785 ;
        RECT 6.41 1.345 6.66 1.785 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.985 1.355 5.68 1.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.85 1.345 6.2 1.675 ;
        RECT 3.645 1.93 6.085 2.1 ;
        RECT 5.85 1.345 6.085 2.1 ;
        RECT 3.645 1.425 3.815 2.1 ;
        RECT 2.805 1.425 3.815 1.625 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 2.265 1.435 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.1168 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.075 0.7 8.255 1.03 ;
        RECT 3.985 0.86 8.255 1.03 ;
        RECT 3.985 0.755 5.965 1.03 ;
        RECT 2.435 1.015 5.605 1.185 ;
        RECT 2.435 1.015 3.815 1.255 ;
        RECT 0.815 1.605 2.635 1.775 ;
        RECT 2.435 1.015 2.635 1.775 ;
        RECT 1.055 0.87 2.605 1.04 ;
        RECT 1.915 0.255 2.105 1.04 ;
        RECT 1.675 1.605 2.005 2.735 ;
        RECT 1.055 0.255 1.245 1.04 ;
        RECT 0.815 1.605 1.145 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.655 -0.085 9.985 1.04 ;
        RECT 8.795 -0.085 9.125 0.7 ;
        RECT 6.135 -0.085 6.465 0.69 ;
        RECT 3.135 -0.085 3.465 0.505 ;
        RECT 2.275 -0.085 2.605 0.7 ;
        RECT 1.415 -0.085 1.745 0.7 ;
        RECT 0.555 -0.085 0.885 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.225 1.945 9.555 3.415 ;
        RECT 8.365 2.295 8.695 3.415 ;
        RECT 7.505 2.295 7.835 3.415 ;
        RECT 6.625 2.295 6.955 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.725 1.605 9.985 3.075 ;
      RECT 8.865 1.605 9.055 3.075 ;
      RECT 8.005 1.955 8.195 3.075 ;
      RECT 7.135 1.955 7.335 3.075 ;
      RECT 2.625 2.77 6.455 3.075 ;
      RECT 6.255 1.955 6.455 3.075 ;
      RECT 6.135 2.27 6.455 3.075 ;
      RECT 2.625 2.285 2.955 3.075 ;
      RECT 6.255 1.955 9.055 2.125 ;
      RECT 8.795 1.605 9.055 2.125 ;
      RECT 8.795 1.605 9.985 1.775 ;
      RECT 8.425 0.87 9.485 1.04 ;
      RECT 9.295 0.255 9.485 1.04 ;
      RECT 8.425 0.255 8.625 1.04 ;
      RECT 6.645 0.255 8.625 0.53 ;
      RECT 0.385 2.905 2.435 3.075 ;
      RECT 2.175 1.945 2.435 3.075 ;
      RECT 1.315 1.945 1.505 3.075 ;
      RECT 0.385 1.815 0.645 3.075 ;
      RECT 3.125 2.27 5.965 2.6 ;
      RECT 3.125 1.795 3.325 2.6 ;
      RECT 2.175 1.945 3.325 2.115 ;
      RECT 3.055 1.795 3.325 2.115 ;
      RECT 2.775 0.675 3.815 0.845 ;
      RECT 3.635 0.255 3.815 0.845 ;
      RECT 2.775 0.505 2.965 0.845 ;
      RECT 3.635 0.255 5.955 0.585 ;
  END
END scs130lp_a221oi_4

MACRO scs130lp_a221oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221oi_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.55 1.385 1.9 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 1 2.755 1.39 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.57 2.755 1.9 ;
        RECT 1.565 1 1.735 1.9 ;
        RECT 1.015 1 1.735 1.33 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.835 1.78 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.945 1.11 3.275 1.78 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5685 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.2 2.04 3.715 3.065 ;
        RECT 3.545 0.265 3.715 3.065 ;
        RECT 1.25 0.65 3.715 0.82 ;
        RECT 3.005 0.265 3.715 0.82 ;
        RECT 1.25 0.265 1.58 0.82 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.07 -0.085 2.4 0.47 ;
        RECT 0.32 -0.085 0.65 0.68 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.32 2.78 1.65 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.67 2.08 3 3.065 ;
      RECT 0.26 2.04 0.59 3.065 ;
      RECT 0.26 2.08 3 2.25 ;
      RECT 2.14 2.43 2.47 3.065 ;
      RECT 0.79 2.43 1.12 3.065 ;
      RECT 0.79 2.43 2.47 2.6 ;
  END
END scs130lp_a221oi_lp

MACRO scs130lp_a221oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a221oi_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.96 1.195 2.245 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.5 0.805 3.205 1.135 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 1.75 3.205 1.965 ;
        RECT 2.555 1.455 3.205 1.965 ;
        RECT 1.5 1.19 1.67 1.965 ;
        RECT 1.34 1.19 1.67 1.36 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.58 1.315 1.93 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.45 1.21 0.805 2.12 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3864 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 0.745 2.245 1.01 ;
        RECT 1.465 0.465 1.795 1.01 ;
        RECT 0.1 2.655 0.865 2.985 ;
        RECT 0.1 0.385 0.515 1.01 ;
        RECT 0.1 0.385 0.27 2.985 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.425 -0.085 2.635 0.585 ;
        RECT 0.735 -0.085 0.945 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.98 2.845 2.31 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.995 2.145 3.205 2.985 ;
      RECT 1.085 2.145 1.295 2.985 ;
      RECT 1.085 2.145 3.205 2.315 ;
      RECT 2.565 2.495 2.775 2.985 ;
      RECT 1.515 2.495 1.725 2.985 ;
      RECT 1.515 2.495 2.775 2.665 ;
  END
END scs130lp_a221oi_m

MACRO scs130lp_a22o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22o_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.795 0.78 3.275 2.19 ;
        RECT 1.385 0.78 3.275 1.015 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 1.185 1.36 1.985 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.185 1.895 1.985 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.185 2.465 1.985 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3105 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.495 0.59 3.075 ;
        RECT 0.085 0.265 0.475 0.595 ;
        RECT 0.085 0.265 0.335 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.41 -0.085 2.74 0.61 ;
        RECT 0.645 -0.085 0.875 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.82 2.445 3.13 3.415 ;
        RECT 0.76 2.495 1.09 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.26 2.905 2.64 3.075 ;
      RECT 2.31 2.445 2.64 3.075 ;
      RECT 1.26 2.505 1.59 3.075 ;
      RECT 1.76 2.155 2.09 2.735 ;
      RECT 0.505 2.155 2.09 2.325 ;
      RECT 0.505 0.775 0.76 2.325 ;
      RECT 0.505 0.775 1.215 0.945 ;
      RECT 1.045 0.28 1.215 0.945 ;
      RECT 1.045 0.28 1.78 0.61 ;
  END
END scs130lp_a22o_0

MACRO scs130lp_a22o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22o_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.33 1.21 2.735 1.56 ;
        RECT 2.45 0.395 2.735 1.56 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.21 3.275 1.56 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.21 2.04 1.48 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.21 1.415 1.48 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 0.255 0.435 1.14 ;
        RECT 0.095 0.255 0.365 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.915 -0.085 3.245 1.04 ;
        RECT 0.605 -0.085 1.345 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.425 2.07 2.765 3.415 ;
        RECT 0.585 1.99 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.935 1.73 3.245 3.075 ;
      RECT 1.045 2.905 2.255 3.075 ;
      RECT 1.975 1.73 2.255 3.075 ;
      RECT 1.045 1.99 1.305 3.075 ;
      RECT 1.975 1.73 3.245 1.9 ;
      RECT 1.475 1.65 1.805 2.735 ;
      RECT 0.605 1.65 1.805 1.82 ;
      RECT 0.605 0.87 0.845 1.82 ;
      RECT 0.605 0.87 2.225 1.04 ;
      RECT 1.895 0.255 2.225 1.04 ;
  END
END scs130lp_a22o_1

MACRO scs130lp_a22o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22o_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.055 1.345 2.245 2.14 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.45 1.345 1.885 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.375 3.745 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.79 1.345 3.205 1.75 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 0.255 0.94 1.065 ;
        RECT 0.605 1.755 0.93 3.075 ;
        RECT 0.57 0.255 0.74 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.595 -0.085 2.925 0.825 ;
        RECT 1.18 -0.085 1.51 0.825 ;
        RECT 0.13 -0.085 0.4 1.105 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.035 2.65 2.365 3.415 ;
        RECT 1.1 1.92 1.43 3.415 ;
        RECT 0.165 2 0.415 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.485 1.93 3.745 3.075 ;
      RECT 2.45 1.93 3.745 2.14 ;
      RECT 2.45 0.995 2.62 2.14 ;
      RECT 0.91 1.245 1.28 1.585 ;
      RECT 1.11 0.995 1.28 1.585 ;
      RECT 1.11 0.995 3.715 1.165 ;
      RECT 3.385 0.255 3.715 1.165 ;
      RECT 2.035 0.255 2.365 1.165 ;
      RECT 2.985 2.31 3.315 3.075 ;
      RECT 1.605 1.92 1.865 3.075 ;
      RECT 1.605 2.31 3.315 2.48 ;
      RECT 1.605 1.92 1.885 2.48 ;
  END
END scs130lp_a22o_2

MACRO scs130lp_a22o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22o_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.31 1.2 6.115 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.77 1.615 6.615 1.785 ;
        RECT 6.285 1.21 6.615 1.785 ;
        RECT 4.77 1.345 5.1 1.785 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.4 1.2 4.02 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.97 1.615 4.56 1.785 ;
        RECT 4.23 1.345 4.56 1.785 ;
        RECT 2.97 1.345 3.23 1.785 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.045 2.46 1.215 ;
        RECT 2.27 0.255 2.46 1.215 ;
        RECT 1.82 1.755 2.05 3.075 ;
        RECT 0.1 1.755 2.05 1.925 ;
        RECT 1.41 0.255 1.59 1.215 ;
        RECT 0.96 1.755 1.15 3.075 ;
        RECT 0.1 0.325 0.425 1.215 ;
        RECT 0.1 0.325 0.345 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 6.335 -0.085 6.625 1.03 ;
        RECT 4.445 -0.085 4.775 0.65 ;
        RECT 2.63 -0.085 2.96 0.65 ;
        RECT 1.77 -0.085 2.1 0.865 ;
        RECT 0.91 -0.085 1.24 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.865 2.295 6.195 3.415 ;
        RECT 4.965 2.295 5.295 3.415 ;
        RECT 2.22 1.815 2.46 3.415 ;
        RECT 1.32 2.095 1.65 3.415 ;
        RECT 0.46 2.095 0.79 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.365 1.955 6.625 3.075 ;
      RECT 5.465 1.955 5.695 3.075 ;
      RECT 2.705 2.905 4.795 3.075 ;
      RECT 4.465 1.955 4.795 3.075 ;
      RECT 3.565 2.305 3.895 3.075 ;
      RECT 2.705 2.305 3.035 3.075 ;
      RECT 4.465 1.955 6.625 2.125 ;
      RECT 5.935 0.255 6.165 1.03 ;
      RECT 5.005 0.255 5.315 0.65 ;
      RECT 5.005 0.255 6.165 0.53 ;
      RECT 4.065 1.955 4.295 2.735 ;
      RECT 3.205 1.955 3.395 2.735 ;
      RECT 2.63 1.955 4.295 2.135 ;
      RECT 2.63 0.82 2.8 2.135 ;
      RECT 0.515 1.385 2.8 1.585 ;
      RECT 2.63 0.82 5.765 1.03 ;
      RECT 5.485 0.7 5.765 1.03 ;
      RECT 3.13 0.255 4.275 0.65 ;
  END
END scs130lp_a22o_4

MACRO scs130lp_a22o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22o_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.795 0.855 2.125 1.185 ;
        RECT 0.415 0.855 2.125 1.025 ;
        RECT 0.125 1.12 0.585 1.79 ;
        RECT 0.415 0.855 0.585 1.79 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.455 1.125 2.785 1.795 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.45 2.275 1.78 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 1.205 1.315 1.875 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.315 2.025 3.725 3.065 ;
        RECT 3.555 0.265 3.725 3.065 ;
        RECT 3.485 1.92 3.725 3.065 ;
        RECT 3.395 0.265 3.725 0.595 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.655 -0.085 2.905 0.595 ;
        RECT 0.67 -0.085 1 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.555 2.325 2.885 3.415 ;
        RECT 0.13 2.025 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.495 1.975 1.825 2.715 ;
      RECT 1.495 1.975 3.135 2.145 ;
      RECT 2.965 0.775 3.135 2.145 ;
      RECT 2.965 0.775 3.375 1.445 ;
      RECT 2.305 0.775 3.375 0.945 ;
      RECT 2.305 0.505 2.475 0.945 ;
      RECT 1.49 0.505 2.475 0.675 ;
      RECT 1.49 0.295 1.82 0.675 ;
      RECT 0.66 2.895 2.355 3.065 ;
      RECT 2.025 2.325 2.355 3.065 ;
      RECT 0.66 2.055 0.99 3.065 ;
  END
END scs130lp_a22o_lp

MACRO scs130lp_a22o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22o_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.615 1.21 3.205 2.49 ;
        RECT 2.445 0.265 2.615 1.38 ;
        RECT 1.535 0.265 2.615 0.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.21 1.325 1.405 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.155 2.245 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.95 2.435 2.12 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.231 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.795 0.64 1.005 ;
        RECT 0.155 2.53 0.55 2.86 ;
        RECT 0.155 0.795 0.325 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.795 -0.085 2.985 0.935 ;
        RECT 0.82 -0.085 1.15 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.84 2.715 3.17 3.415 ;
        RECT 0.73 2.675 1.06 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.3 2.895 2.66 3.065 ;
      RECT 2.45 2.675 2.66 3.065 ;
      RECT 1.3 2.675 1.63 3.065 ;
      RECT 1.845 2.325 2.175 2.715 ;
      RECT 0.765 2.325 2.175 2.495 ;
      RECT 0.765 1.585 0.935 2.495 ;
      RECT 0.505 1.585 0.935 2.255 ;
      RECT 0.505 1.585 1.795 1.755 ;
      RECT 1.625 0.645 1.795 1.755 ;
      RECT 1.625 0.645 1.93 0.975 ;
  END
END scs130lp_a22o_m

MACRO scs130lp_a22oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22oi_0 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 0.39 1.775 1.485 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 0.765 2.315 1.485 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 0.765 1.295 1.485 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.8 0.375 1.835 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3556 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 0.265 1.295 0.595 ;
        RECT 0.625 1.665 0.945 2.685 ;
        RECT 0.545 0.265 0.715 1.835 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.945 -0.085 2.275 0.595 ;
        RECT 0.125 -0.085 0.375 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.54 2.005 1.81 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.185 2.855 1.37 3.025 ;
      RECT 1.115 1.665 1.37 3.025 ;
      RECT 0.185 2.005 0.455 3.025 ;
      RECT 1.98 1.665 2.27 2.685 ;
      RECT 1.115 1.665 2.27 1.835 ;
  END
END scs130lp_a22oi_0

MACRO scs130lp_a22oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22oi_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.18 1.845 1.75 ;
        RECT 1.585 1.1 1.845 1.75 ;
        RECT 1.585 0.365 1.81 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 1.21 2.795 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.21 1.35 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.535 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.693 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.705 1.92 2.245 2.13 ;
        RECT 0.705 0.86 1.415 1.04 ;
        RECT 1.205 0.325 1.415 1.04 ;
        RECT 0.705 1.92 1.045 2.735 ;
        RECT 0.705 0.86 0.875 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.17 -0.085 2.5 0.995 ;
        RECT 0.285 -0.085 0.535 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.63 2.64 2.3 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.47 1.92 2.73 3.075 ;
      RECT 0.285 2.905 1.46 3.075 ;
      RECT 1.215 2.3 1.46 3.075 ;
      RECT 0.285 1.92 0.535 3.075 ;
      RECT 1.215 2.3 2.73 2.47 ;
      RECT 2.415 1.92 2.73 2.47 ;
  END
END scs130lp_a22oi_1

MACRO scs130lp_a22oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22oi_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.95 2.375 2.12 ;
        RECT 2.125 1.345 2.375 2.12 ;
        RECT 0.625 1.345 0.885 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.345 1.915 1.78 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.985 1.345 4.555 1.75 ;
        RECT 2.905 1.925 4.165 2.095 ;
        RECT 3.985 1.345 4.165 2.095 ;
        RECT 2.905 1.345 3.155 2.095 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.365 1.345 3.815 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6044 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.55 1.005 4.68 1.175 ;
        RECT 4.4 0.255 4.68 1.175 ;
        RECT 3.92 2.265 4.24 2.595 ;
        RECT 2.55 2.265 4.24 2.435 ;
        RECT 0.44 0.995 2.74 1.165 ;
        RECT 2.55 0.255 2.735 2.435 ;
        RECT 2.41 0.255 2.74 1.165 ;
        RECT 0.44 0.255 0.69 1.165 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.49 -0.085 3.82 0.495 ;
        RECT 1.38 -0.085 1.71 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 1.71 2.945 2.41 3.415 ;
        RECT 1.71 2.63 2.04 3.415 ;
        RECT 0.75 2.63 1.08 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.59 2.765 4.68 3.075 ;
      RECT 4.41 1.99 4.68 3.075 ;
      RECT 1.28 2.29 1.54 3.075 ;
      RECT 0.205 2.29 0.535 3.075 ;
      RECT 2.21 2.605 3.725 2.775 ;
      RECT 2.21 2.29 2.38 2.775 ;
      RECT 0.205 2.29 2.38 2.46 ;
      RECT 0.205 1.855 0.455 3.075 ;
      RECT 2.98 0.665 4.23 0.835 ;
      RECT 3.99 0.505 4.23 0.835 ;
      RECT 2.98 0.255 3.32 0.835 ;
      RECT 0.87 0.655 2.22 0.825 ;
      RECT 1.89 0.265 2.22 0.825 ;
      RECT 0.87 0.265 1.2 0.825 ;
  END
END scs130lp_a22oi_2

MACRO scs130lp_a22oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22oi_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.88 1.21 6.58 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.75 1.425 8.005 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.775 1.355 4.645 1.525 ;
        RECT 2.985 1.21 4.645 1.525 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.12 1.21 2.245 1.525 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 0.815 5.845 1.04 ;
        RECT 5.645 0.695 5.845 1.04 ;
        RECT 3.495 1.705 3.825 2.735 ;
        RECT 0.835 1.705 3.825 1.875 ;
        RECT 2.555 1.705 2.885 2.735 ;
        RECT 2.425 0.595 2.815 1.145 ;
        RECT 2.425 0.595 2.595 1.875 ;
        RECT 1.695 1.705 2.025 2.735 ;
        RECT 0.835 1.705 1.165 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.305 -0.085 7.635 0.895 ;
        RECT 6.445 -0.085 6.775 0.605 ;
        RECT 1.565 -0.085 1.895 0.7 ;
        RECT 0.705 -0.085 1.035 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.085 2.27 7.415 3.415 ;
        RECT 6.225 2.27 6.555 3.415 ;
        RECT 5.32 2.095 5.65 3.415 ;
        RECT 4.46 2.095 4.79 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.855 1.065 8.065 1.255 ;
      RECT 7.805 0.255 8.065 1.255 ;
      RECT 6.855 0.775 7.135 1.255 ;
      RECT 6.945 0.255 7.135 1.255 ;
      RECT 6.015 0.775 7.135 1.04 ;
      RECT 6.015 0.275 6.275 1.04 ;
      RECT 4.295 0.275 6.275 0.525 ;
      RECT 7.585 1.93 7.845 3.075 ;
      RECT 6.725 1.93 6.915 3.075 ;
      RECT 5.82 1.93 6.055 3.075 ;
      RECT 4.96 1.755 5.15 3.075 ;
      RECT 0.405 2.905 4.29 3.075 ;
      RECT 3.995 1.755 4.29 3.075 ;
      RECT 3.055 2.045 3.325 3.075 ;
      RECT 2.195 2.045 2.385 3.075 ;
      RECT 1.335 2.045 1.525 3.075 ;
      RECT 0.405 1.825 0.665 3.075 ;
      RECT 5.82 1.93 7.845 2.1 ;
      RECT 5.82 1.755 6.045 3.075 ;
      RECT 3.995 1.755 6.045 1.925 ;
      RECT 0.275 0.87 2.245 1.04 ;
      RECT 2.065 0.255 2.245 1.04 ;
      RECT 1.205 0.315 1.395 1.04 ;
      RECT 0.275 0.315 0.535 1.04 ;
      RECT 2.995 0.255 4.045 0.635 ;
      RECT 2.065 0.255 4.045 0.425 ;
  END
END scs130lp_a22oi_4

MACRO scs130lp_a22oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22oi_lp 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.575 1.075 1.965 1.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.33 0.855 2.755 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 1.075 1.395 1.745 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 1.075 0.855 1.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4438 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.725 1.55 0.895 ;
        RECT 1.22 0.265 1.55 0.895 ;
        RECT 0.83 1.925 1.16 2.715 ;
        RECT 0.125 1.925 1.16 2.095 ;
        RECT 0.125 0.725 0.345 2.095 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.33 -0.085 2.66 0.675 ;
        RECT 0.4 -0.085 0.73 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.89 2.275 2.22 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.43 1.925 2.76 3.065 ;
      RECT 0.3 2.895 1.69 3.065 ;
      RECT 1.36 1.925 1.69 3.065 ;
      RECT 0.3 2.275 0.63 3.065 ;
      RECT 1.36 1.925 2.76 2.095 ;
  END
END scs130lp_a22oi_lp

MACRO scs130lp_a22oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a22oi_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.505 0.47 1.765 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 0.84 2.245 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.96 0.84 1.285 2.12 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.49 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2835 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.61 0.33 1.27 0.66 ;
        RECT 0.685 2.32 1.015 2.71 ;
        RECT 0.61 0.33 0.78 2.49 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.945 -0.085 2.275 0.485 ;
        RECT 0.24 -0.085 0.43 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.545 2.67 1.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.175 2.89 1.365 3.06 ;
      RECT 1.195 2.32 1.365 3.06 ;
      RECT 0.175 2.67 0.505 3.06 ;
      RECT 2.055 2.32 2.245 2.79 ;
      RECT 1.195 2.32 2.245 2.49 ;
  END
END scs130lp_a22oi_m

MACRO scs130lp_a2bb2o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2o_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.53 0.78 0.935 1.76 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.145 1.655 1.75 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.42 0.4 3.755 2.195 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.76 0.78 3.25 2.195 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2935 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.28 0.595 0.61 ;
        RECT 0.085 2.43 0.445 3.075 ;
        RECT 0.085 0.28 0.335 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.98 -0.085 3.25 0.61 ;
        RECT 1.66 -0.085 1.99 0.61 ;
        RECT 0.765 -0.085 1.025 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.02 2.755 3.285 3.415 ;
        RECT 0.615 2.43 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.455 2.415 3.745 3.05 ;
      RECT 2.59 2.415 2.825 3.05 ;
      RECT 2.59 2.415 3.745 2.585 ;
      RECT 1.14 2.88 2.42 3.05 ;
      RECT 2.185 2.075 2.42 3.05 ;
      RECT 1.14 1.93 1.31 3.05 ;
      RECT 0.505 1.93 1.31 2.26 ;
      RECT 2.325 0.28 2.495 2.245 ;
      RECT 2.16 0.28 2.495 0.61 ;
      RECT 1.48 2.43 2.005 2.71 ;
      RECT 1.835 0.78 2.005 2.71 ;
      RECT 1.835 1.235 2.155 1.905 ;
      RECT 1.195 0.78 2.005 0.975 ;
      RECT 1.195 0.28 1.465 0.975 ;
  END
END scs130lp_a2bb2o_0

MACRO scs130lp_a2bb2o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2o_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 0.37 1.295 2.155 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.015 1.925 1.525 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 0.84 3.755 2.225 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.915 0.28 3.215 2.225 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.815 0.565 3.075 ;
        RECT 0.105 0.255 0.505 1.095 ;
        RECT 0.105 0.255 0.285 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.385 -0.085 3.655 0.61 ;
        RECT 1.89 -0.085 2.22 0.495 ;
        RECT 0.675 -0.085 0.935 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.93 2.735 3.26 3.415 ;
        RECT 0.735 2.665 1.065 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.43 2.395 3.69 3.02 ;
      RECT 2.535 2.395 2.76 3.02 ;
      RECT 2.535 2.395 3.69 2.565 ;
      RECT 2.07 2.325 2.365 3.02 ;
      RECT 2.17 2.055 2.365 3.02 ;
      RECT 0.755 2.325 2.365 2.495 ;
      RECT 0.755 1.345 0.925 2.495 ;
      RECT 2.17 2.055 2.735 2.225 ;
      RECT 2.565 0.28 2.735 2.225 ;
      RECT 0.455 1.345 0.925 1.645 ;
      RECT 2.45 0.28 2.735 0.675 ;
      RECT 1.78 1.705 1.99 2.145 ;
      RECT 1.78 1.705 2.385 1.875 ;
      RECT 2.11 1.005 2.385 1.875 ;
      RECT 2.11 0.665 2.28 1.875 ;
      RECT 1.465 0.665 2.28 0.835 ;
      RECT 1.465 0.28 1.715 0.835 ;
  END
END scs130lp_a2bb2o_1

MACRO scs130lp_a2bb2o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2o_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.21 2.87 2.13 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.96 1.21 2.375 1.435 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.185 0.395 2.215 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.565 1.185 1.02 2.215 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.38 1.85 3.74 3.075 ;
        RECT 3.57 0.255 3.74 3.075 ;
        RECT 3.37 0.255 3.74 1.095 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.91 -0.085 4.12 1.095 ;
        RECT 2.94 -0.085 3.13 0.885 ;
        RECT 1.61 -0.085 1.94 0.68 ;
        RECT 0.275 -0.085 0.605 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.91 1.815 4.12 3.415 ;
        RECT 2.88 2.64 3.21 3.415 ;
        RECT 0.545 2.725 0.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.46 2.3 1.755 3.055 ;
      RECT 1.46 2.3 3.21 2.47 ;
      RECT 3.04 1.34 3.21 2.47 ;
      RECT 1.46 2.045 1.695 3.055 ;
      RECT 1.19 2.045 1.695 2.215 ;
      RECT 1.19 0.685 1.36 2.215 ;
      RECT 3.04 1.34 3.4 1.67 ;
      RECT 1.065 0.685 1.36 1.015 ;
      RECT 1.945 1.685 2.275 2.13 ;
      RECT 1.53 1.685 2.275 1.855 ;
      RECT 1.53 0.86 1.79 1.855 ;
      RECT 1.53 0.86 2.625 1.03 ;
      RECT 2.415 0.7 2.625 1.03 ;
      RECT 0.095 2.385 0.365 3.075 ;
      RECT 1.055 2.385 1.29 3.065 ;
      RECT 0.095 2.385 1.29 2.555 ;
  END
END scs130lp_a2bb2o_2

MACRO scs130lp_a2bb2o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2o_4 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.475 1.065 5.04 1.515 ;
        RECT 3.245 1.065 5.04 1.235 ;
        RECT 3.245 1.065 3.575 1.435 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 1.415 4.295 1.75 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.405 1.97 1.645 ;
        RECT 0.545 1.95 1.635 2.12 ;
        RECT 1.465 1.405 1.635 2.12 ;
        RECT 0.545 1.345 0.715 2.12 ;
        RECT 0.24 1.345 0.715 1.645 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 1.405 1.295 1.78 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1886 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.55 1.755 7.045 1.925 ;
        RECT 6.875 1.065 7.045 1.925 ;
        RECT 5.475 1.065 7.045 1.235 ;
        RECT 6.41 1.755 6.63 3.075 ;
        RECT 6.375 0.255 6.565 1.235 ;
        RECT 5.55 1.755 5.74 3.075 ;
        RECT 5.475 0.255 5.705 1.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 6.735 -0.085 7.065 0.895 ;
        RECT 5.875 -0.085 6.205 0.865 ;
        RECT 5.025 -0.085 5.305 0.885 ;
        RECT 4.015 -0.085 4.345 0.555 ;
        RECT 2.735 -0.085 3.405 0.555 ;
        RECT 1.905 -0.085 2.185 0.895 ;
        RECT 0.115 -0.085 0.4 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.8 2.095 7.1 3.415 ;
        RECT 5.91 2.095 6.24 3.415 ;
        RECT 5.02 2.65 5.35 3.415 ;
        RECT 3.255 2.65 3.585 3.415 ;
        RECT 1.425 2.63 1.755 3.415 ;
        RECT 0.545 2.63 0.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.345 1.065 2.565 2.735 ;
      RECT 2.365 0.255 2.565 2.735 ;
      RECT 3.235 2.31 5.38 2.48 ;
      RECT 5.21 1.405 5.38 2.48 ;
      RECT 3.235 2.1 3.405 2.48 ;
      RECT 2.345 2.1 3.405 2.27 ;
      RECT 5.21 1.405 6.695 1.585 ;
      RECT 1.02 1.065 2.565 1.235 ;
      RECT 1.02 0.595 1.235 1.235 ;
      RECT 3.575 1.93 4.445 2.14 ;
      RECT 2.755 1.76 3.745 1.93 ;
      RECT 2.755 0.725 2.925 1.93 ;
      RECT 2.755 0.725 4.855 0.895 ;
      RECT 4.525 0.255 4.855 0.895 ;
      RECT 3.575 0.255 3.835 0.895 ;
      RECT 1.935 2.905 3.065 3.075 ;
      RECT 2.735 2.44 3.065 3.075 ;
      RECT 1.045 2.29 1.255 3.075 ;
      RECT 0.095 1.815 0.375 3.075 ;
      RECT 1.935 1.815 2.175 3.075 ;
      RECT 0.095 2.29 2.175 2.46 ;
      RECT 0.57 0.255 0.85 1.095 ;
      RECT 1.405 0.255 1.735 0.895 ;
      RECT 0.57 0.255 1.735 0.425 ;
      RECT 3.755 2.67 4.85 3 ;
  END
END scs130lp_a2bb2o_4

MACRO scs130lp_a2bb2o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2o_lp 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 1.18 3.89 2.15 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 1.11 5.155 1.78 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.17 1.345 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.17 0.835 1.84 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.68 1.92 3.235 2.15 ;
        RECT 2.68 1.92 3.055 2.325 ;
        RECT 2.68 0.35 2.85 2.325 ;
        RECT 2.465 0.35 2.85 0.81 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.835 -0.085 5.165 0.81 ;
        RECT 3.255 -0.085 3.585 0.81 ;
        RECT 1.115 -0.085 1.445 0.64 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 3.335 2.835 3.665 3.415 ;
        RECT 0.725 2.37 1.055 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.265 2.025 4.765 3.065 ;
      RECT 1.765 2.495 4.765 2.665 ;
      RECT 4.095 0.35 4.265 2.665 ;
      RECT 1.765 1.17 1.935 2.665 ;
      RECT 1.6 1.17 1.935 1.84 ;
      RECT 4.045 0.35 4.375 0.81 ;
      RECT 2.115 0.99 2.445 2.325 ;
      RECT 2.115 0.99 2.5 1.66 ;
      RECT 1.905 0.265 2.235 0.99 ;
      RECT 0.295 0.82 2.285 0.99 ;
      RECT 0.295 0.265 0.625 0.99 ;
      RECT 1.255 2.02 1.585 3.06 ;
      RECT 0.195 2.02 0.525 3.06 ;
      RECT 0.195 2.02 1.585 2.19 ;
  END
END scs130lp_a2bb2o_lp

MACRO scs130lp_a2bb2o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2o_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.21 1.765 1.405 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.95 1.765 2.49 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 1.21 3.685 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.47 2.855 1.825 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.145 2.655 0.48 2.985 ;
        RECT 0.145 0.47 0.475 0.875 ;
        RECT 0.145 0.47 0.325 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.27 -0.085 3.6 0.875 ;
        RECT 0.655 0.86 1.865 1.03 ;
        RECT 1.675 0.7 1.865 1.03 ;
        RECT 0.655 -0.085 0.865 1.03 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.82 2.355 3.15 3.415 ;
        RECT 0.66 2.845 0.99 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.36 2.005 3.57 2.455 ;
      RECT 2.43 2.005 2.64 2.455 ;
      RECT 2.43 2.005 3.57 2.175 ;
      RECT 2 1.6 2.215 2.435 ;
      RECT 2.045 0.795 2.215 2.435 ;
      RECT 0.505 1.6 0.675 2.395 ;
      RECT 0.505 1.6 2.215 1.77 ;
      RECT 2.045 0.795 2.375 1.38 ;
      RECT 1.105 0.265 1.435 0.68 ;
      RECT 1.105 0.265 2.25 0.435 ;
      RECT 1.45 2.735 2.315 3.065 ;
  END
END scs130lp_a2bb2o_m

MACRO scs130lp_a2bb2oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2oi_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.455 1.84 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 0.78 1.365 1.435 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.865 0.78 3.275 1.475 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.055 0.78 2.55 1.475 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2872 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.715 0.275 2.28 0.61 ;
        RECT 1.57 1.915 1.935 2.95 ;
        RECT 1.57 0.78 1.885 2.95 ;
        RECT 1.715 0.275 1.885 2.95 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.91 -0.085 3.24 0.61 ;
        RECT 1 -0.085 1.545 0.61 ;
        RECT 0.095 -0.085 0.385 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.505 1.985 2.835 3.415 ;
        RECT 0.095 2.115 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.015 1.645 3.265 2.595 ;
      RECT 2.105 1.645 2.335 2.595 ;
      RECT 2.105 1.645 3.265 1.815 ;
      RECT 0.885 1.645 1.215 2.795 ;
      RECT 0.625 1.645 1.4 2.155 ;
      RECT 0.625 0.28 0.83 2.155 ;
      RECT 0.555 0.28 0.83 0.61 ;
  END
END scs130lp_a2bb2oi_0

MACRO scs130lp_a2bb2oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2oi_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.805 1.75 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.975 1.185 1.385 1.515 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.915 1.21 3.275 1.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.2 2.405 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5691 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.45 2.035 2.745 2.205 ;
        RECT 2.575 0.86 2.745 2.205 ;
        RECT 1.95 0.86 2.745 1.03 ;
        RECT 1.95 0.255 2.15 1.03 ;
        RECT 1.45 2.035 1.775 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.925 -0.085 3.195 1.04 ;
        RECT 0.97 -0.085 1.78 0.675 ;
        RECT 0.11 -0.085 0.44 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.38 2.715 2.71 3.415 ;
        RECT 0.11 1.92 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.88 2.375 3.195 3.075 ;
      RECT 2.915 1.93 3.195 3.075 ;
      RECT 1.945 2.375 2.21 3.075 ;
      RECT 1.945 2.375 3.195 2.545 ;
      RECT 0.93 1.92 1.26 3.075 ;
      RECT 0.975 1.695 1.26 3.075 ;
      RECT 0.975 1.695 1.735 1.865 ;
      RECT 1.555 0.845 1.735 1.865 ;
      RECT 1.555 1.2 1.895 1.515 ;
      RECT 0.61 0.845 1.735 1.015 ;
      RECT 0.61 0.255 0.8 1.015 ;
  END
END scs130lp_a2bb2oi_1

MACRO scs130lp_a2bb2oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2oi_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 1.415 3.955 1.875 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.175 1.21 5.675 1.75 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.425 2.015 1.655 ;
        RECT 0.55 1.92 1.88 2.12 ;
        RECT 1.595 1.425 1.88 2.12 ;
        RECT 0.55 1.375 0.73 2.12 ;
        RECT 0.235 1.375 0.73 1.625 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.91 1.425 1.425 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8232 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.42 1.805 2.75 2.735 ;
        RECT 2.5 0.285 2.75 2.735 ;
        RECT 0.97 1.075 2.75 1.245 ;
        RECT 2.49 0.285 2.75 1.245 ;
        RECT 0.97 0.605 1.3 1.245 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 5.175 -0.085 5.505 1.04 ;
        RECT 4.315 -0.085 4.645 0.895 ;
        RECT 2.92 -0.085 3.785 0.895 ;
        RECT 1.99 -0.085 2.32 0.895 ;
        RECT 0.11 -0.085 0.405 1.185 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 3.885 2.385 4.215 3.415 ;
        RECT 1.49 2.63 1.82 3.415 ;
        RECT 0.54 2.63 0.87 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.385 2.905 5.505 3.075 ;
      RECT 5.175 1.92 5.505 3.075 ;
      RECT 3.455 2.045 3.715 3.075 ;
      RECT 4.385 2.045 4.615 3.075 ;
      RECT 3.455 2.045 4.615 2.215 ;
      RECT 4.785 1.705 5.005 2.735 ;
      RECT 4.135 1.705 5.005 1.875 ;
      RECT 4.135 1.075 4.305 1.875 ;
      RECT 3.085 1.075 3.335 1.605 ;
      RECT 3.085 1.075 4.995 1.245 ;
      RECT 4.825 0.305 4.995 1.245 ;
      RECT 3.955 0.305 4.145 1.245 ;
      RECT 2.05 2.905 3.18 3.075 ;
      RECT 2.92 1.825 3.18 3.075 ;
      RECT 1.04 2.29 1.24 3.075 ;
      RECT 0.11 1.815 0.37 3.075 ;
      RECT 2.05 1.825 2.25 3.075 ;
      RECT 0.11 2.29 2.25 2.46 ;
      RECT 0.11 1.815 0.38 2.46 ;
      RECT 0.575 0.265 0.8 1.185 ;
      RECT 1.47 0.265 1.82 0.905 ;
      RECT 0.575 0.265 1.82 0.435 ;
  END
END scs130lp_a2bb2oi_2

MACRO scs130lp_a2bb2oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2oi_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.22 1.405 8.04 1.755 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.21 1.345 9.56 1.525 ;
        RECT 8.21 1.21 8.965 1.525 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.635 1.665 3.825 1.835 ;
        RECT 3.505 1.2 3.825 1.835 ;
        RECT 1.635 1.35 1.805 1.835 ;
        RECT 0.295 1.35 1.805 1.555 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.985 1.315 3.335 1.485 ;
        RECT 2.04 1.2 3.335 1.485 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.355 1.045 5.7 1.38 ;
        RECT 5.215 1.89 5.545 2.735 ;
        RECT 5.215 0.255 5.405 1.215 ;
        RECT 3.995 1.89 5.545 2.085 ;
        RECT 4.345 1.045 5.7 1.215 ;
        RECT 3.995 1.885 4.77 2.085 ;
        RECT 4.355 1.885 4.685 2.735 ;
        RECT 4.345 0.255 4.545 1.215 ;
        RECT 2.05 0.755 4.545 1.03 ;
        RECT 4.31 0.255 4.545 1.03 ;
        RECT 3.995 0.755 4.165 2.085 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.535 -0.085 9.865 0.835 ;
        RECT 8.675 -0.085 9.005 0.7 ;
        RECT 7.295 -0.085 8.135 0.7 ;
        RECT 7.295 -0.085 7.625 0.87 ;
        RECT 6.435 -0.085 6.765 0.895 ;
        RECT 5.575 -0.085 5.905 0.875 ;
        RECT 4.715 -0.085 5.045 0.865 ;
        RECT 3.81 -0.085 4.14 0.585 ;
        RECT 1.19 -0.085 1.52 0.84 ;
        RECT 0.33 -0.085 0.62 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 7.455 2.27 7.785 3.415 ;
        RECT 6.595 2.27 6.925 3.415 ;
        RECT 3.415 2.585 3.745 3.415 ;
        RECT 2.475 2.355 2.805 3.415 ;
        RECT 1.615 2.355 1.945 3.415 ;
        RECT 0.755 2.065 1.085 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.215 1.695 9.475 2.735 ;
      RECT 8.34 1.695 8.615 2.735 ;
      RECT 8.34 1.695 9.935 1.875 ;
      RECT 9.73 1.005 9.935 1.875 ;
      RECT 4.94 1.55 6.05 1.72 ;
      RECT 5.88 1.065 6.05 1.72 ;
      RECT 4.335 1.385 5.185 1.715 ;
      RECT 5.88 1.065 8.04 1.235 ;
      RECT 9.165 1.005 9.935 1.175 ;
      RECT 6.935 1.04 8.04 1.235 ;
      RECT 6.075 0.255 6.265 1.235 ;
      RECT 7.87 0.87 9.365 1.04 ;
      RECT 6.935 0.255 7.125 1.235 ;
      RECT 9.175 0.255 9.365 1.175 ;
      RECT 8.305 0.255 8.505 1.04 ;
      RECT 7.955 2.905 9.935 3.075 ;
      RECT 9.645 2.045 9.935 3.075 ;
      RECT 7.095 1.93 7.285 3.075 ;
      RECT 6.165 1.93 6.425 3.075 ;
      RECT 8.785 2.045 9.045 3.075 ;
      RECT 7.955 1.93 8.17 3.075 ;
      RECT 6.165 1.93 8.17 2.1 ;
      RECT 3.915 2.905 5.975 3.075 ;
      RECT 5.715 1.89 5.975 3.075 ;
      RECT 2.975 2.015 3.175 3.075 ;
      RECT 2.115 2.015 2.305 3.075 ;
      RECT 1.255 1.725 1.445 3.075 ;
      RECT 0.325 1.725 0.585 3.075 ;
      RECT 4.855 2.255 5.045 3.075 ;
      RECT 3.915 2.255 4.185 3.075 ;
      RECT 3.845 2.255 4.185 2.425 ;
      RECT 2.975 2.245 3.905 2.415 ;
      RECT 2.975 2.015 3.715 2.415 ;
      RECT 1.255 2.015 3.715 2.185 ;
      RECT 1.255 1.725 1.465 2.185 ;
      RECT 0.325 1.725 1.465 1.895 ;
      RECT 0.79 1.01 1.87 1.18 ;
      RECT 1.69 0.255 1.87 1.18 ;
      RECT 0.79 0.255 1.02 1.18 ;
      RECT 1.69 0.255 3.64 0.585 ;
  END
END scs130lp_a2bb2oi_4

MACRO scs130lp_a2bb2oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2oi_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.475 1.11 4.195 1.78 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 0.775 2.845 1.105 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.81 0.835 1.14 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.45 1.315 1.78 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3976 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.705 1.635 2.035 3.065 ;
        RECT 1.085 0.265 1.795 0.675 ;
        RECT 1.495 1.635 2.035 1.805 ;
        RECT 1.495 0.265 1.665 1.805 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.595 -0.085 3.925 0.675 ;
        RECT 2.005 -0.085 2.335 0.675 ;
        RECT 0.395 -0.085 0.725 0.63 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.88 2.025 4.21 3.415 ;
        RECT 0.645 2.335 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.26 2.895 3.68 3.065 ;
      RECT 3.35 2.025 3.68 3.065 ;
      RECT 2.26 1.675 2.59 3.065 ;
      RECT 2.79 1.285 3.12 2.715 ;
      RECT 1.845 1.285 3.195 1.455 ;
      RECT 3.025 0.265 3.195 1.455 ;
      RECT 1.845 1.125 2.175 1.455 ;
      RECT 2.805 0.265 3.195 0.595 ;
      RECT 1.175 1.985 1.505 3.065 ;
      RECT 0.115 1.985 0.445 3.065 ;
      RECT 0.115 1.985 1.505 2.155 ;
  END
END scs130lp_a2bb2oi_lp

MACRO scs130lp_a2bb2oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a2bb2oi_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.47 0.355 2.49 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 0.895 2.86 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 0.765 3.205 1.435 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.195 0.765 2.725 1.435 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.845 0.375 2.21 0.585 ;
        RECT 1.595 1.405 2.015 1.575 ;
        RECT 1.845 0.375 2.015 1.575 ;
        RECT 1.595 1.405 1.83 2.245 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.78 -0.085 3.11 0.485 ;
        RECT 1.475 -0.085 1.665 0.545 ;
        RECT 0.535 -0.085 0.865 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.42 2.105 2.75 3.415 ;
        RECT 0.125 2.755 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.93 1.755 3.12 2.245 ;
      RECT 2.05 1.755 2.24 2.245 ;
      RECT 2.05 1.755 3.12 1.925 ;
      RECT 1.075 2.695 1.695 3.025 ;
      RECT 1.075 0.33 1.265 3.025 ;
      RECT 1.045 0.33 1.265 0.66 ;
  END
END scs130lp_a2bb2oi_m

MACRO scs130lp_a311o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311o_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 0.37 2.29 1.865 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 0.37 1.83 1.865 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.98 0.77 1.365 1.86 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.46 1.08 2.83 1.865 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.37 1.08 3.755 2.22 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2937 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.41 0.565 3.075 ;
        RECT 0.085 0.285 0.565 1.39 ;
        RECT 0.085 0.285 0.26 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.895 -0.085 3.205 0.57 ;
        RECT 0.735 -0.085 1.065 0.6 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.635 2.74 2.165 3.415 ;
        RECT 0.735 2.41 0.965 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.02 2.39 3.455 3.075 ;
      RECT 3.02 0.74 3.2 3.075 ;
      RECT 0.43 2.035 3.2 2.23 ;
      RECT 3 0.74 3.2 2.23 ;
      RECT 0.43 1.56 0.69 2.23 ;
      RECT 2.48 0.74 3.645 0.91 ;
      RECT 3.375 0.285 3.645 0.91 ;
      RECT 2.48 0.285 2.725 0.91 ;
      RECT 1.135 2.4 1.465 3.075 ;
      RECT 2.335 2.4 2.665 3.02 ;
      RECT 1.135 2.4 2.665 2.57 ;
  END
END scs130lp_a311o_0

MACRO scs130lp_a311o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311o_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.195 2.365 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.195 1.905 1.525 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 1.195 1.365 1.525 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.535 1.195 3.215 1.525 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.195 3.755 1.525 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.035 0.67 3.075 ;
        RECT 0.085 0.255 0.355 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.88 -0.085 3.21 0.685 ;
        RECT 0.525 -0.085 1.24 0.685 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.7 2.375 2.38 3.415 ;
        RECT 0.84 2.035 1.1 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.38 1.695 3.71 3.075 ;
      RECT 0.605 1.695 3.71 1.865 ;
      RECT 0.605 0.855 0.84 1.865 ;
      RECT 0.525 0.855 0.84 1.515 ;
      RECT 0.525 0.855 3.71 1.025 ;
      RECT 3.38 0.255 3.71 1.025 ;
      RECT 2.325 0.255 2.655 1.025 ;
      RECT 2.55 2.035 2.88 3.075 ;
      RECT 1.27 2.035 1.53 3.075 ;
      RECT 1.27 2.035 2.88 2.205 ;
  END
END scs130lp_a311o_1

MACRO scs130lp_a311o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311o_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.185 2.835 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 1.185 2.335 1.525 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.445 1.185 1.825 1.525 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.185 3.695 1.525 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.865 1.185 4.235 1.525 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.85 0.905 3.075 ;
        RECT 0.635 0.255 0.81 3.075 ;
        RECT 0.58 0.255 0.81 1.535 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.25 -0.085 3.58 0.675 ;
        RECT 0.98 -0.085 1.65 0.675 ;
        RECT 0.12 -0.085 0.41 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.26 2.385 2.59 3.415 ;
        RECT 1.15 2.045 1.48 3.415 ;
        RECT 0.195 1.815 0.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.73 1.695 4.06 3.075 ;
      RECT 1.075 1.695 4.06 1.875 ;
      RECT 1.075 0.845 1.245 1.875 ;
      RECT 0.985 0.845 1.245 1.515 ;
      RECT 0.985 0.845 4.06 1.015 ;
      RECT 3.75 0.255 4.06 1.015 ;
      RECT 2.705 0.255 3.035 1.015 ;
      RECT 2.83 2.045 3.16 3.065 ;
      RECT 1.68 2.045 2.01 3.065 ;
      RECT 1.68 2.045 3.16 2.215 ;
  END
END scs130lp_a311o_2

MACRO scs130lp_a311o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311o_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.315 1.21 7.595 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.775 1.345 6.375 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.895 1.415 5.605 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.97 1.415 1.865 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.43 1.75 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4304 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.06 1.405 4.725 1.75 ;
        RECT 2.99 1.75 4.395 2.015 ;
        RECT 4.06 1.025 4.23 2.015 ;
        RECT 2.375 1.025 4.23 1.195 ;
        RECT 3.23 0.255 3.42 1.195 ;
        RECT 2.375 0.255 2.56 1.195 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 4.79 -0.085 5.12 0.845 ;
        RECT 3.59 -0.085 4.26 0.855 ;
        RECT 2.73 -0.085 3.06 0.855 ;
        RECT 1.86 -0.085 2.19 0.905 ;
        RECT 0.975 -0.085 1.305 0.905 ;
        RECT 0.1 -0.085 0.43 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.245 1.92 7.575 3.415 ;
        RECT 6.345 2.6 6.675 3.415 ;
        RECT 5.45 2.6 5.78 3.415 ;
        RECT 4.59 2.865 4.92 3.415 ;
        RECT 3.48 2.865 3.81 3.415 ;
        RECT 2.465 2.865 2.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.415 0.255 6.645 1.175 ;
      RECT 7.315 0.255 7.575 1.04 ;
      RECT 5.45 0.255 5.745 0.835 ;
      RECT 5.45 0.255 7.575 0.425 ;
      RECT 0.6 0.255 0.79 2.735 ;
      RECT 2.64 2.185 4.735 2.355 ;
      RECT 4.565 1.92 4.735 2.355 ;
      RECT 2.64 1.365 2.81 2.355 ;
      RECT 4.565 1.92 6.715 2.09 ;
      RECT 6.545 1.345 6.715 2.09 ;
      RECT 6.545 1.345 7.145 1.645 ;
      RECT 6.815 0.595 7.145 1.645 ;
      RECT 2.035 1.365 2.81 1.585 ;
      RECT 2.035 1.365 3.865 1.535 ;
      RECT 2.035 1.075 2.205 1.585 ;
      RECT 0.6 1.075 2.205 1.245 ;
      RECT 1.475 0.255 1.69 1.245 ;
      RECT 0.6 0.255 0.805 1.245 ;
      RECT 6.845 2.26 7.075 3.075 ;
      RECT 6.885 1.815 7.075 3.075 ;
      RECT 5.95 2.26 6.16 3.075 ;
      RECT 5.09 2.26 5.28 3.075 ;
      RECT 1.46 1.92 1.69 2.735 ;
      RECT 2.29 2.525 5.28 2.695 ;
      RECT 5.02 2.26 5.28 2.695 ;
      RECT 2.29 1.92 2.46 2.695 ;
      RECT 5.02 2.26 7.075 2.43 ;
      RECT 1.46 1.92 2.46 2.09 ;
      RECT 4.43 1.065 5.38 1.235 ;
      RECT 5.915 0.595 6.245 1.175 ;
      RECT 5.21 1.005 6.245 1.175 ;
      RECT 4.43 0.255 4.62 1.235 ;
      RECT 0.1 2.905 2.12 3.075 ;
      RECT 1.86 2.26 2.12 3.075 ;
      RECT 0.96 1.92 1.29 3.075 ;
      RECT 0.1 1.92 0.43 3.075 ;
  END
END scs130lp_a311o_4

MACRO scs130lp_a311o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311o_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.2 2.755 1.87 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.2 1.865 1.87 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 1.2 1.325 1.87 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 1.24 3.265 2.89 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 1.2 3.835 1.87 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.265 0.835 0.67 ;
        RECT 0.105 2.05 0.53 3.065 ;
        RECT 0.105 0.265 0.275 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.015 -0.085 3.345 0.67 ;
        RECT 1.015 -0.085 1.345 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 1.79 2.4 2.12 3.415 ;
        RECT 0.73 2.05 1.06 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.73 2.05 4.185 3.065 ;
      RECT 4.015 0.85 4.185 3.065 ;
      RECT 0.455 0.85 0.785 1.52 ;
      RECT 0.455 0.85 4.185 1.02 ;
      RECT 3.805 0.265 4.135 1.02 ;
      RECT 2.225 0.265 2.555 1.02 ;
      RECT 2.425 2.05 2.755 3.065 ;
      RECT 1.26 2.05 1.59 3.065 ;
      RECT 1.26 2.05 2.755 2.22 ;
  END
END scs130lp_a311o_lp

MACRO scs130lp_a311o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311o_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.74 1.58 2.245 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.47 1.53 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 0.91 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.01 2.43 1.38 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.21 3.205 1.75 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.35 0.425 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.245 -0.085 2.575 0.47 ;
        RECT 0.605 -0.085 0.935 0.49 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.465 2.28 1.795 3.415 ;
        RECT 0.605 2.125 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.975 2.855 2.78 3.025 ;
      RECT 2.61 0.65 2.78 3.025 ;
      RECT 2.61 2.055 3.095 2.265 ;
      RECT 1.855 0.65 3.035 0.82 ;
      RECT 2.825 0.35 3.035 0.82 ;
      RECT 1.855 0.35 2.065 0.82 ;
      RECT 2.035 1.93 2.245 2.325 ;
      RECT 1.015 1.93 1.225 2.325 ;
      RECT 1.015 1.93 2.245 2.1 ;
  END
END scs130lp_a311o_m

MACRO scs130lp_a311oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311oi_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.485 1.155 1.82 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 0.4 1.315 1.825 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 0.78 0.84 1.835 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.075 2.32 2.66 ;
        RECT 1.99 1.075 2.32 1.86 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.49 1.13 2.86 2.175 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4111 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.495 2.345 3.275 3.025 ;
        RECT 3.03 0.28 3.275 3.025 ;
        RECT 1.595 0.735 3.275 0.905 ;
        RECT 2.855 0.28 3.275 0.905 ;
        RECT 1.595 0.28 1.92 0.905 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.09 -0.085 2.685 0.565 ;
        RECT 0.105 -0.085 0.775 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.23 2.345 1.5 3.415 ;
        RECT 0.335 2.355 0.63 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.67 2.005 1.895 3.025 ;
      RECT 0.8 2.005 1.06 3.025 ;
      RECT 0.8 2.005 1.895 2.175 ;
  END
END scs130lp_a311oi_0

MACRO scs130lp_a311oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311oi_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.185 1.905 1.52 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 1.185 1.375 1.52 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.19 0.89 1.52 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.185 2.475 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.985 1.185 3.235 1.515 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9093 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.97 1.705 3.265 3.075 ;
        RECT 1.035 0.84 3.265 1.015 ;
        RECT 2.935 0.255 3.265 1.015 ;
        RECT 2.645 1.705 3.265 1.875 ;
        RECT 2.645 0.84 2.815 1.875 ;
        RECT 1.035 0.255 2.245 1.015 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.425 -0.085 2.755 0.67 ;
        RECT 0.45 -0.085 0.78 1.02 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.46 2.03 1.79 3.415 ;
        RECT 0.45 1.815 0.78 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.075 1.69 2.405 3.075 ;
      RECT 0.95 1.69 1.235 3.075 ;
      RECT 0.95 1.69 2.405 1.86 ;
  END
END scs130lp_a311oi_1

MACRO scs130lp_a311oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311oi_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.29 1.425 3.685 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.94 1.415 2.735 1.75 ;
        RECT 1.385 1.415 2.735 1.585 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.415 1.105 1.585 ;
        RECT 0.155 1.415 0.55 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.9 1.425 4.23 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.4 1.425 5.675 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3524 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.085 5.665 1.255 ;
        RECT 5.385 0.305 5.665 1.255 ;
        RECT 4.92 1.92 5.195 2.735 ;
        RECT 1.975 1.92 5.195 2.12 ;
        RECT 4.525 0.305 4.715 1.255 ;
        RECT 3.665 0.305 3.855 1.255 ;
        RECT 2.905 1.085 3.075 2.12 ;
        RECT 2.655 0.595 2.995 1.245 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.885 -0.085 5.215 0.915 ;
        RECT 4.025 -0.085 4.355 0.915 ;
        RECT 0.65 -0.085 0.98 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 3.035 2.63 3.365 3.415 ;
        RECT 2.06 2.63 2.39 3.415 ;
        RECT 1.08 2.095 1.41 3.415 ;
        RECT 0.22 1.92 0.55 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.595 2.905 5.645 3.075 ;
      RECT 5.365 1.92 5.645 3.075 ;
      RECT 3.595 2.8 4.75 3.075 ;
      RECT 4.49 2.29 4.75 3.075 ;
      RECT 2.605 2.29 2.865 3.075 ;
      RECT 1.58 2.29 1.84 3.075 ;
      RECT 0.72 1.755 0.9 3.075 ;
      RECT 4.025 2.29 4.32 2.63 ;
      RECT 1.58 2.29 4.32 2.46 ;
      RECT 1.58 1.755 1.77 3.075 ;
      RECT 0.72 1.755 1.77 1.925 ;
      RECT 1.51 0.255 1.84 0.905 ;
      RECT 3.165 0.255 3.495 0.895 ;
      RECT 1.51 0.255 3.495 0.425 ;
      RECT 0.22 1.075 2.35 1.245 ;
      RECT 2.01 0.595 2.35 1.245 ;
      RECT 1.15 0.325 1.34 1.245 ;
      RECT 0.22 0.325 0.48 1.245 ;
  END
END scs130lp_a311oi_2

MACRO scs130lp_a311oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311oi_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.345 1.21 5.695 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.01 1.21 3.81 1.435 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 1.84 1.435 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.865 1.21 7.7 1.435 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.91 1.21 9.995 1.435 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.3352 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.995 0.87 9.655 1.04 ;
        RECT 9.395 0.255 9.655 1.04 ;
        RECT 9.035 1.605 9.265 2.735 ;
        RECT 3.995 1.605 9.265 1.775 ;
        RECT 8.535 0.255 8.725 1.04 ;
        RECT 8.175 1.605 8.365 2.735 ;
        RECT 7.62 0.255 7.865 1.04 ;
        RECT 6.715 0.255 6.95 1.04 ;
        RECT 5.805 0.255 6.045 1.04 ;
        RECT 4.95 0.655 5.21 1.04 ;
        RECT 3.995 0.655 4.355 1.04 ;
        RECT 3.995 0.655 4.175 1.775 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.895 -0.085 9.225 0.7 ;
        RECT 8.035 -0.085 8.365 0.7 ;
        RECT 7.12 -0.085 7.45 0.7 ;
        RECT 6.215 -0.085 6.545 0.7 ;
        RECT 1.385 -0.085 1.715 0.7 ;
        RECT 0.525 -0.085 0.855 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 5.435 2.285 5.765 3.415 ;
        RECT 4.575 2.285 4.905 3.415 ;
        RECT 3.66 2.285 3.99 3.415 ;
        RECT 2.745 1.945 3.075 3.415 ;
        RECT 1.885 1.945 2.215 3.415 ;
        RECT 1.025 1.945 1.355 3.415 ;
        RECT 0.165 1.815 0.495 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.955 2.905 9.725 3.075 ;
      RECT 9.435 1.815 9.725 3.075 ;
      RECT 8.535 1.945 8.865 3.075 ;
      RECT 7.675 1.945 8.005 3.075 ;
      RECT 6.815 2.285 7.145 3.075 ;
      RECT 5.955 2.285 6.285 3.075 ;
      RECT 5.075 1.945 5.265 3.075 ;
      RECT 4.16 1.945 4.405 3.075 ;
      RECT 3.245 1.605 3.49 3.075 ;
      RECT 2.385 1.605 2.575 3.075 ;
      RECT 1.525 1.605 1.715 3.075 ;
      RECT 0.665 1.605 0.855 3.075 ;
      RECT 7.315 1.945 7.505 2.735 ;
      RECT 6.455 1.945 6.645 2.735 ;
      RECT 3.245 1.945 7.505 2.115 ;
      RECT 3.245 1.605 3.505 2.115 ;
      RECT 0.665 1.605 3.505 1.775 ;
      RECT 5.38 0.255 5.635 0.7 ;
      RECT 4.525 0.255 4.78 0.7 ;
      RECT 3.135 0.255 3.4 0.7 ;
      RECT 2.285 0.255 2.54 0.7 ;
      RECT 3.135 0.255 5.635 0.485 ;
      RECT 2.285 0.255 5.635 0.445 ;
      RECT 0.095 0.87 3.825 1.04 ;
      RECT 3.57 0.665 3.825 1.04 ;
      RECT 2.71 0.665 2.965 1.04 ;
      RECT 1.885 0.255 2.115 1.04 ;
      RECT 1.025 0.255 1.215 1.04 ;
      RECT 0.095 0.255 0.355 1.04 ;
  END
END scs130lp_a311oi_4

MACRO scs130lp_a311oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311oi_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.81 0.58 1.14 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.51 1.21 1.84 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.42 1.17 1.795 1.84 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 1.17 2.32 1.84 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.345 2.89 1.78 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5223 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.785 2.025 3.24 3.065 ;
        RECT 3.07 0.81 3.24 3.065 ;
        RECT 3.005 0.81 3.24 1.04 ;
        RECT 0.76 0.82 3.24 0.99 ;
        RECT 2.125 0.265 2.455 0.99 ;
        RECT 0.76 0.46 0.93 0.99 ;
        RECT 0.125 0.46 0.93 0.63 ;
        RECT 0.125 0.265 0.455 0.63 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.915 -0.085 3.245 0.63 ;
        RECT 1.335 -0.085 1.665 0.64 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.175 2.37 1.505 3.415 ;
        RECT 0.115 2.025 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.725 2.02 2.055 3.065 ;
      RECT 0.645 2.02 0.975 3.065 ;
      RECT 0.645 2.02 2.055 2.19 ;
  END
END scs130lp_a311oi_lp

MACRO scs130lp_a311oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a311oi_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.775 2.205 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 0.47 1.285 2.12 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 0.47 0.805 2.86 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.315 2.12 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 2.855 2.49 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3423 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.645 2.67 3.205 3 ;
        RECT 3.035 0.365 3.205 3 ;
        RECT 1.75 0.685 3.205 0.855 ;
        RECT 2.63 0.365 3.205 0.855 ;
        RECT 1.75 0.365 1.94 0.855 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.12 -0.085 2.45 0.505 ;
        RECT 0.155 -0.085 0.345 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.42 2.805 1.61 3.415 ;
        RECT 0.155 2.785 0.345 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.99 2.455 1.2 2.965 ;
      RECT 1.79 2.455 2.12 2.925 ;
      RECT 0.99 2.455 2.12 2.625 ;
  END
END scs130lp_a311oi_m

MACRO scs130lp_a31o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31o_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.01 0.795 2.39 1.51 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.575 0.795 1.84 1.51 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 1.01 1.36 1.52 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.995 0.795 3.275 1.84 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2893 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.395 0.74 3.075 ;
        RECT 0.085 0.27 0.555 0.5 ;
        RECT 0.085 0.27 0.34 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.775 -0.085 3.105 0.625 ;
        RECT 0.735 -0.085 1.065 0.5 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.775 2.395 2.025 3.415 ;
        RECT 0.91 2.395 1.17 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.625 2.395 2.925 3.075 ;
      RECT 2.625 1.705 2.825 3.075 ;
      RECT 0.51 1.705 2.825 1.875 ;
      RECT 0.51 0.67 0.76 1.875 ;
      RECT 0.51 0.67 1.405 0.84 ;
      RECT 1.235 0.295 1.405 0.84 ;
      RECT 1.235 0.295 2.605 0.625 ;
      RECT 2.195 2.055 2.455 3.075 ;
      RECT 1.34 2.055 1.605 3.075 ;
      RECT 1.34 2.055 2.455 2.225 ;
  END
END scs130lp_a31o_0

MACRO scs130lp_a31o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31o_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.055 1.21 2.375 1.54 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.555 1.21 1.885 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.975 1.21 1.345 1.54 ;
        RECT 1.095 1.21 1.285 2.86 ;
        RECT 0.975 1.21 1.285 1.645 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.21 2.925 1.54 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.695 0.405 3.075 ;
        RECT 0.085 0.255 0.345 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.79 -0.085 3.12 0.7 ;
        RECT 0.525 -0.085 1.22 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.865 2.05 2.195 3.415 ;
        RECT 0.625 1.815 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.83 1.815 3.12 3.075 ;
      RECT 3.095 0.87 3.265 1.985 ;
      RECT 0.515 0.87 0.765 1.515 ;
      RECT 0.515 0.87 3.265 1.04 ;
      RECT 2.29 0.255 2.62 1.04 ;
      RECT 2.365 1.71 2.66 3.075 ;
      RECT 1.455 1.71 1.695 3.075 ;
      RECT 1.455 1.71 2.66 1.88 ;
  END
END scs130lp_a31o_1

MACRO scs130lp_a31o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31o_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.485 1.195 3.215 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.985 1.195 2.315 1.525 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 1.195 1.815 1.525 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.195 3.755 1.525 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 2.045 1.05 3.065 ;
        RECT 0.635 0.255 0.81 3.065 ;
        RECT 0.62 0.255 0.81 1.125 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.19 -0.085 3.52 1.025 ;
        RECT 0.98 -0.085 1.65 0.685 ;
        RECT 0.12 -0.085 0.45 1.1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.225 2.445 2.555 3.415 ;
        RECT 1.22 2.045 1.55 3.415 ;
        RECT 0.205 1.825 0.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.26 1.705 3.52 3.075 ;
      RECT 0.985 1.705 3.52 1.875 ;
      RECT 0.985 1.195 1.345 1.875 ;
      RECT 1.175 0.855 1.345 1.875 ;
      RECT 1.175 0.855 3.02 1.025 ;
      RECT 2.69 0.255 3.02 1.025 ;
      RECT 1.72 2.045 2.015 3.075 ;
      RECT 2.76 2.045 3.09 3.065 ;
      RECT 1.72 2.045 3.09 2.225 ;
  END
END scs130lp_a31o_2

MACRO scs130lp_a31o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31o_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.915 1.415 6.565 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.955 1.415 5.605 1.76 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.515 1.415 4.645 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.425 1.76 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5932 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.405 1.93 3.575 2.26 ;
        RECT 1.025 0.975 2.9 1.185 ;
        RECT 1.405 0.975 1.69 2.26 ;
        RECT 1.025 0.975 1.69 1.76 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 4.105 -0.085 4.305 0.545 ;
        RECT 3.095 -0.085 3.425 0.465 ;
        RECT 2.045 -0.085 2.375 0.465 ;
        RECT 0.955 -0.085 1.285 0.465 ;
        RECT 0.095 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 6.295 1.93 6.625 3.415 ;
        RECT 5.435 2.27 5.765 3.415 ;
        RECT 4.555 2.27 4.885 3.415 ;
        RECT 3.675 2.78 4.005 3.415 ;
        RECT 2.815 2.78 3.145 3.415 ;
        RECT 1.955 2.78 2.285 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.365 0.275 6.625 1.195 ;
      RECT 5.515 0.275 5.695 0.645 ;
      RECT 4.575 0.275 5.695 0.555 ;
      RECT 4.575 0.275 6.625 0.445 ;
      RECT 0.595 0.635 0.855 2.735 ;
      RECT 1.89 1.355 3.25 1.645 ;
      RECT 3.08 0.635 3.25 1.645 ;
      RECT 3.08 1.075 6.195 1.245 ;
      RECT 5.865 0.615 6.195 1.245 ;
      RECT 0.595 0.635 3.25 0.805 ;
      RECT 0.595 0.255 0.785 2.735 ;
      RECT 5.935 1.93 6.125 3.075 ;
      RECT 5.055 1.93 5.265 3.075 ;
      RECT 4.175 1.93 4.385 3.075 ;
      RECT 0.095 2.905 1.285 3.075 ;
      RECT 1.025 2.44 1.285 3.075 ;
      RECT 0.095 1.93 0.425 3.075 ;
      RECT 1.025 2.44 4.385 2.61 ;
      RECT 4.105 1.93 4.385 2.61 ;
      RECT 1.025 1.93 1.235 3.075 ;
      RECT 4.105 1.93 6.125 2.1 ;
      RECT 3.605 0.725 5.335 0.905 ;
      RECT 3.605 0.345 3.935 0.905 ;
  END
END scs130lp_a31o_4

MACRO scs130lp_a31o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31o_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.165 1.315 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 0.44 1.855 1.495 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.165 2.395 1.495 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.445 1.165 0.805 1.495 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.87 2.025 3.27 3.065 ;
        RECT 3.1 0.265 3.27 3.065 ;
        RECT 2.915 0.265 3.27 0.72 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.125 -0.085 2.455 0.72 ;
        RECT 0.125 -0.085 0.455 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.34 2.025 2.67 3.415 ;
        RECT 1.28 2.375 1.61 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.095 1.675 0.55 3.065 ;
      RECT 0.095 1.675 2.92 1.845 ;
      RECT 2.605 1.175 2.92 1.845 ;
      RECT 0.095 0.815 0.265 3.065 ;
      RECT 0.095 0.815 1.245 0.985 ;
      RECT 0.915 0.265 1.245 0.985 ;
      RECT 1.81 2.025 2.14 3.065 ;
      RECT 0.75 2.025 1.08 3.065 ;
      RECT 0.75 2.025 2.14 2.195 ;
  END
END scs130lp_a31o_lp

MACRO scs130lp_a31o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31o_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.3 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.59 1.21 1.765 2.12 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.05 1.21 1.285 2.49 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 2.87 2.49 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 1.71 0.735 2.87 ;
        RECT 0.155 0.35 0.725 0.68 ;
        RECT 0.155 1.71 0.735 1.88 ;
        RECT 0.155 0.35 0.325 1.88 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.595 -0.085 2.805 0.64 ;
        RECT 0.905 -0.085 1.235 0.58 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.835 2.67 2.025 3.415 ;
        RECT 0.915 2.73 1.245 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.715 2.67 2.905 3 ;
      RECT 2.715 2.67 3.22 2.84 ;
      RECT 3.05 0.86 3.22 2.84 ;
      RECT 0.51 0.86 0.68 1.53 ;
      RECT 0.51 0.86 3.22 1.03 ;
      RECT 2.165 0.44 2.375 1.03 ;
      RECT 1.425 2.67 1.635 3 ;
      RECT 1.465 2.32 1.635 3 ;
      RECT 2.205 2.67 2.535 2.88 ;
      RECT 2.205 2.32 2.375 2.88 ;
      RECT 1.465 2.32 2.375 2.49 ;
  END
END scs130lp_a31o_m

MACRO scs130lp_a31oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31oi_0 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.095 0.785 1.505 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.39 0.925 1.825 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.765 0.455 1.82 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 0.84 2.315 1.78 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.346 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.845 1.95 2.315 3.025 ;
        RECT 1.675 0.28 1.845 2.175 ;
        RECT 1.375 0.28 1.845 0.615 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 2.015 -0.085 2.295 0.61 ;
        RECT 0.125 -0.085 0.455 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.99 1.995 1.25 2.735 ;
        RECT 0.095 1.995 1.25 2.165 ;
        RECT 0.095 1.995 0.39 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.56 2.905 1.675 3.075 ;
      RECT 1.42 2.345 1.675 3.075 ;
      RECT 0.56 2.345 0.82 3.075 ;
  END
END scs130lp_a31oi_0

MACRO scs130lp_a31oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31oi_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 1.185 1.845 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 0.75 1.345 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.545 1.78 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 1.185 2.795 1.515 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7623 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.25 1.685 2.795 3.075 ;
        RECT 0.715 1.685 2.795 1.855 ;
        RECT 1.635 0.255 2.01 1.015 ;
        RECT 0.715 0.255 2.01 0.53 ;
        RECT 0.715 0.255 0.885 1.855 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.18 -0.085 2.51 1.015 ;
        RECT 0.3 -0.085 0.545 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.24 2.365 1.57 3.415 ;
        RECT 0.3 1.95 0.56 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.75 2.025 2.08 3.065 ;
      RECT 0.73 2.025 1.06 3.065 ;
      RECT 0.73 2.025 2.08 2.195 ;
  END
END scs130lp_a31oi_1

MACRO scs130lp_a31oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31oi_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.96 1.425 3.335 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.21 1.635 1.545 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 1.21 0.455 1.545 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 1.425 4.715 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0374 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.335 1.085 4.465 1.255 ;
        RECT 4.205 0.325 4.465 1.255 ;
        RECT 3.705 1.95 4.035 2.735 ;
        RECT 2.335 1.95 4.035 2.13 ;
        RECT 3.345 0.325 3.535 1.255 ;
        RECT 2.335 1.085 2.79 2.13 ;
        RECT 2.335 0.605 2.675 2.13 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.705 -0.085 4.035 0.915 ;
        RECT 0.525 -0.085 0.855 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 2.325 2.64 3.175 3.415 ;
        RECT 1.43 2.055 1.76 3.415 ;
        RECT 0.525 2.055 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.345 2.905 4.465 3.075 ;
      RECT 4.205 1.92 4.465 3.075 ;
      RECT 1.93 1.715 2.155 3.075 ;
      RECT 1.025 1.715 1.26 3.075 ;
      RECT 0.095 1.715 0.355 3.075 ;
      RECT 3.345 2.3 3.535 3.075 ;
      RECT 1.93 2.3 3.535 2.47 ;
      RECT 1.93 1.715 2.165 2.47 ;
      RECT 0.095 1.715 2.165 1.885 ;
      RECT 2.845 0.255 3.175 0.915 ;
      RECT 1.425 0.255 1.645 0.7 ;
      RECT 1.425 0.255 3.175 0.435 ;
      RECT 1.815 0.605 2.145 1.205 ;
      RECT 0.095 0.87 2.145 1.04 ;
      RECT 1.025 0.335 1.255 1.04 ;
      RECT 0.095 0.335 0.345 1.04 ;
  END
END scs130lp_a31oi_2

MACRO scs130lp_a31oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31oi_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.875 1.425 6.565 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.93 1.425 4.165 1.76 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.425 2.725 1.76 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.75 1.425 8.06 1.78 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8564 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.355 1.075 8.065 1.255 ;
        RECT 7.815 0.305 8.065 1.255 ;
        RECT 7.235 1.95 7.565 2.735 ;
        RECT 4.355 1.95 7.565 2.12 ;
        RECT 6.945 0.285 7.135 1.255 ;
        RECT 6.375 1.95 6.705 2.735 ;
        RECT 4.355 1.05 6.275 1.255 ;
        RECT 6.075 0.285 6.275 1.255 ;
        RECT 4.355 0.84 5.485 1.255 ;
        RECT 5.155 0.595 5.485 1.255 ;
        RECT 4.355 0.84 4.705 2.12 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.305 -0.085 7.635 0.905 ;
        RECT 6.445 -0.085 6.775 0.905 ;
        RECT 1.385 -0.085 1.715 0.915 ;
        RECT 0.525 -0.085 0.855 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 5.435 2.63 5.765 3.415 ;
        RECT 4.575 2.63 4.905 3.415 ;
        RECT 3.175 2.64 4.015 3.415 ;
        RECT 3.175 2.27 3.845 3.415 ;
        RECT 2.315 2.27 2.645 3.415 ;
        RECT 1.455 2.27 1.785 3.415 ;
        RECT 0.595 2.27 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.935 2.905 7.995 3.075 ;
      RECT 7.745 1.95 7.995 3.075 ;
      RECT 5.075 2.29 5.265 3.075 ;
      RECT 4.185 2.29 4.405 3.075 ;
      RECT 2.815 1.93 3.005 3.075 ;
      RECT 1.955 1.93 2.145 3.075 ;
      RECT 1.095 1.93 1.285 3.075 ;
      RECT 0.165 1.93 0.425 3.075 ;
      RECT 6.875 2.29 7.065 3.075 ;
      RECT 5.935 2.29 6.205 3.075 ;
      RECT 4.015 1.93 4.185 2.47 ;
      RECT 4.015 2.29 6.205 2.46 ;
      RECT 0.165 1.93 4.185 2.1 ;
      RECT 3.265 0.255 3.595 0.915 ;
      RECT 2.245 0.255 2.575 0.915 ;
      RECT 5.655 0.255 5.855 0.88 ;
      RECT 4.725 0.255 4.985 0.67 ;
      RECT 2.245 0.255 5.855 0.425 ;
      RECT 0.095 1.085 4.105 1.255 ;
      RECT 3.775 0.595 4.105 1.255 ;
      RECT 2.755 0.595 3.085 1.255 ;
      RECT 1.885 0.325 2.075 1.255 ;
      RECT 1.025 0.325 1.215 1.255 ;
      RECT 0.095 0.325 0.345 1.255 ;
  END
END scs130lp_a31oi_4

MACRO scs130lp_a31oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31oi_lp 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.505 1.12 1.835 1.79 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.935 0.44 1.315 1.79 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.695 1.78 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.12 2.405 1.79 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.3 2.025 2.755 3.065 ;
        RECT 2.585 0.77 2.755 3.065 ;
        RECT 1.63 0.77 2.755 0.94 ;
        RECT 1.63 0.265 1.96 0.94 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.42 -0.085 2.75 0.59 ;
        RECT 0.42 -0.085 0.75 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.2 2.32 1.53 3.415 ;
        RECT 0.14 2.025 0.47 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.77 1.97 2.1 3.065 ;
      RECT 0.67 1.97 1 3.065 ;
      RECT 0.67 1.97 2.1 2.14 ;
  END
END scs130lp_a31oi_lp

MACRO scs130lp_a31oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a31oi_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.47 1.765 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 0.47 1.285 2.12 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.49 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.305 1.88 ;
        RECT 2.075 1.21 2.245 2.12 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3507 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.17 2.48 2.725 2.81 ;
        RECT 2.555 0.84 2.725 2.81 ;
        RECT 1.97 0.84 2.725 1.01 ;
        RECT 1.97 0.52 2.18 1.01 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.36 -0.085 2.69 0.66 ;
        RECT 0.49 -0.085 0.82 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.25 2.69 1.58 3.415 ;
        RECT 0.39 2.67 0.72 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.76 2.34 1.95 2.79 ;
      RECT 0.9 2.34 1.07 2.79 ;
      RECT 0.9 2.34 1.95 2.51 ;
  END
END scs130lp_a31oi_m

MACRO scs130lp_a32o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32o_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.02 0.78 2.375 1.51 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.015 1.85 1.685 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.965 1.015 1.35 1.745 ;
        RECT 0.965 1.015 1.305 1.86 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 0.78 2.915 1.51 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.425 0.78 3.755 1.85 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.125 0.755 2.935 ;
        RECT 0.085 0.255 0.355 0.585 ;
        RECT 0.085 0.255 0.335 2.935 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.425 -0.085 3.675 0.61 ;
        RECT 0.525 -0.085 1.25 0.505 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.865 2.205 2.195 3.415 ;
        RECT 0.925 2.125 1.205 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.365 2.895 3.6 3.065 ;
      RECT 3.32 2.125 3.6 3.065 ;
      RECT 2.365 1.865 2.65 3.065 ;
      RECT 1.375 2.03 1.695 2.805 ;
      RECT 1.475 1.865 2.65 2.035 ;
      RECT 2.82 1.785 3.15 2.725 ;
      RECT 3.085 0.28 3.255 1.955 ;
      RECT 0.505 0.675 0.755 1.955 ;
      RECT 0.505 0.675 1.85 0.845 ;
      RECT 1.595 0.28 1.85 0.845 ;
      RECT 1.595 0.28 3.255 0.61 ;
  END
END scs130lp_a32o_0

MACRO scs130lp_a32o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32o_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.195 2.365 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.195 1.875 1.525 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.195 1.35 1.525 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.195 3.25 1.515 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.42 1.21 3.755 1.75 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.85 0.545 3.075 ;
        RECT 0.095 0.255 0.345 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.38 -0.085 3.71 1.04 ;
        RECT 0.545 -0.085 1.195 0.685 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.65 2.385 2.38 3.415 ;
        RECT 0.72 2.105 1.05 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.55 2.905 3.71 3.075 ;
      RECT 3.42 1.93 3.71 3.075 ;
      RECT 1.22 2.045 1.48 3.065 ;
      RECT 2.55 2.045 2.75 3.075 ;
      RECT 1.22 2.045 2.75 2.215 ;
      RECT 2.92 1.705 3.25 2.735 ;
      RECT 0.715 1.705 3.25 1.875 ;
      RECT 0.715 0.855 0.885 1.875 ;
      RECT 0.515 0.855 0.885 1.515 ;
      RECT 0.515 0.855 2.92 1.025 ;
      RECT 2.24 0.255 2.92 1.025 ;
  END
END scs130lp_a32o_1

MACRO scs130lp_a32o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32o_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 0.36 3.255 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.425 0.36 4.165 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.345 1.21 4.715 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.185 2.735 2.575 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.345 2.015 1.76 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.903 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.165 1.775 1.415 3.075 ;
        RECT 0.155 1.775 1.415 1.945 ;
        RECT 0.155 1.065 1.075 1.235 ;
        RECT 0.885 0.255 1.075 1.235 ;
        RECT 0.155 1.065 0.875 1.945 ;
        RECT 0.155 1.065 0.495 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.335 -0.085 4.59 1.04 ;
        RECT 1.245 -0.085 2.035 0.835 ;
        RECT 0.385 -0.085 0.715 0.895 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.21 1.92 4.54 3.415 ;
        RECT 3.3 2.105 3.63 3.415 ;
        RECT 0.665 2.115 0.995 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.8 1.755 4.04 3.075 ;
      RECT 1.685 2.905 3.13 3.075 ;
      RECT 2.905 1.755 3.13 3.075 ;
      RECT 2.565 2.745 3.13 3.075 ;
      RECT 1.685 1.93 2.015 3.075 ;
      RECT 2.905 1.755 4.04 1.925 ;
      RECT 2.185 1.005 2.375 2.735 ;
      RECT 1.085 1.405 1.415 1.605 ;
      RECT 1.245 1.005 1.415 1.605 ;
      RECT 1.245 1.005 2.375 1.175 ;
      RECT 2.205 0.255 2.865 1.005 ;
  END
END scs130lp_a32o_2

MACRO scs130lp_a32o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32o_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.18 1.435 6.085 1.75 ;
        RECT 5.425 1.355 6.085 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.455 1.415 4.205 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.54 1.425 3.245 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.615 1.425 7.045 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.355 1.425 8.005 1.75 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.74 1.755 1.97 3.075 ;
        RECT 0.1 1.045 1.82 1.215 ;
        RECT 1.56 0.255 1.82 1.215 ;
        RECT 0.1 1.755 1.97 1.925 ;
        RECT 0.88 1.755 1.07 3.075 ;
        RECT 0.7 0.255 0.89 1.215 ;
        RECT 0.1 1.045 0.335 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.29 -0.085 7.62 0.905 ;
        RECT 3.03 -0.085 3.24 0.565 ;
        RECT 2.01 -0.085 2.34 0.905 ;
        RECT 1.06 -0.085 1.39 0.875 ;
        RECT 0.2 -0.085 0.53 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 5.27 2.26 5.6 3.415 ;
        RECT 4.41 2.26 4.74 3.415 ;
        RECT 2.96 2.26 3.29 3.415 ;
        RECT 2.14 1.815 2.37 3.415 ;
        RECT 1.24 2.095 1.57 3.415 ;
        RECT 0.38 2.095 0.71 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.93 1.075 8.05 1.245 ;
      RECT 7.79 0.255 8.05 1.245 ;
      RECT 6.93 0.255 7.12 1.245 ;
      RECT 6 0.255 6.26 0.835 ;
      RECT 6 0.255 7.12 0.425 ;
      RECT 5.77 2.905 8.04 3.075 ;
      RECT 7.78 1.92 8.04 3.075 ;
      RECT 4.91 1.92 5.1 3.075 ;
      RECT 3.865 1.92 4.24 3.075 ;
      RECT 2.54 1.92 2.79 3.075 ;
      RECT 6.775 2.27 7.105 3.075 ;
      RECT 5.77 1.92 6.085 3.075 ;
      RECT 2.54 1.92 6.085 2.09 ;
      RECT 7.28 1.92 7.61 2.735 ;
      RECT 6.255 1.92 6.535 2.735 ;
      RECT 6.255 1.92 7.61 2.1 ;
      RECT 6.255 1.005 6.435 2.735 ;
      RECT 0.505 1.385 2.195 1.585 ;
      RECT 2.025 1.075 2.195 1.585 ;
      RECT 4.35 1.095 5.255 1.265 ;
      RECT 2.025 1.075 4.52 1.245 ;
      RECT 6.43 0.595 6.76 1.175 ;
      RECT 5.065 1.005 6.76 1.175 ;
      RECT 5.065 0.615 5.31 1.175 ;
      RECT 4.69 0.255 4.895 0.925 ;
      RECT 3.76 0.685 4.895 0.895 ;
      RECT 5.48 0.255 5.81 0.835 ;
      RECT 4.69 0.255 5.81 0.445 ;
      RECT 2.53 0.735 3.58 0.905 ;
      RECT 3.41 0.255 3.58 0.905 ;
      RECT 2.53 0.255 2.86 0.905 ;
      RECT 3.41 0.255 4.52 0.515 ;
  END
END scs130lp_a32o_4

MACRO scs130lp_a32o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32o_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.235 1.825 1.905 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 0.81 2.395 1.905 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.925 1.55 3.255 1.88 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.925 1.235 1.315 1.905 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.235 0.685 1.905 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4425 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.865 0.44 4.205 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 2.925 -0.085 3.175 1.02 ;
        RECT 0.23 -0.085 0.56 1.055 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.925 2.075 3.255 3.415 ;
        RECT 1.72 2.785 2.05 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.66 2.085 0.99 2.715 ;
      RECT 0.66 2.085 2.745 2.255 ;
      RECT 2.575 0.46 2.745 2.255 ;
      RECT 2.575 1.2 3.685 1.37 ;
      RECT 3.355 0.265 3.685 1.37 ;
      RECT 1.19 0.46 1.52 1.055 ;
      RECT 1.19 0.46 2.745 0.63 ;
      RECT 2.33 2.435 2.66 3.065 ;
      RECT 0.13 2.895 1.52 3.065 ;
      RECT 1.19 2.435 1.52 3.065 ;
      RECT 0.13 2.085 0.46 3.065 ;
      RECT 1.19 2.435 2.66 2.605 ;
  END
END scs130lp_a32o_lp

MACRO scs130lp_a32o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32o_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.97 0.765 2.245 1.095 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.35 0.47 1.765 1.015 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 1.14 1.015 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 2.69 3.205 2.965 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 0.84 3.205 1.75 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.231 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.905 0.425 2.235 ;
        RECT 0.155 0.33 0.395 0.66 ;
        RECT 0.155 0.33 0.325 2.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.915 -0.085 3.245 0.485 ;
        RECT 0.575 -0.085 0.905 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 0.605 2.335 1.815 2.505 ;
        RECT 1.625 2.035 1.815 2.505 ;
        RECT 0.605 1.945 0.935 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.035 2.335 3.125 2.505 ;
      RECT 2.915 2.035 3.125 2.505 ;
      RECT 2.035 1.685 2.225 2.505 ;
      RECT 1.115 1.685 1.445 2.155 ;
      RECT 1.115 1.685 2.225 1.855 ;
      RECT 2.405 1.945 2.735 2.155 ;
      RECT 2.565 0.375 2.735 2.155 ;
      RECT 0.505 1.335 0.675 1.665 ;
      RECT 0.505 1.335 2.735 1.505 ;
      RECT 2.125 0.375 2.735 0.585 ;
  END
END scs130lp_a32o_m

MACRO scs130lp_a32oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32oi_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 0.385 1.85 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.02 0.385 2.415 1.445 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.66 0.78 3.275 1.795 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 0.775 1.36 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.455 1.795 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3556 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.265 1.36 0.595 ;
        RECT 0.625 0.265 0.855 2.645 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.75 -0.085 3.08 0.61 ;
        RECT 0.245 -0.085 0.455 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.66 1.965 2.965 3.415 ;
        RECT 1.47 1.965 2.075 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.145 2.815 1.3 2.985 ;
      RECT 1.025 1.615 1.3 2.985 ;
      RECT 0.145 1.965 0.455 2.985 ;
      RECT 2.245 1.615 2.49 2.645 ;
      RECT 1.025 1.615 2.49 1.795 ;
  END
END scs130lp_a32oi_0

MACRO scs130lp_a32oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32oi_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 0.37 1.835 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 0.37 2.35 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.52 1.21 3.275 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.02 1.21 1.365 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.51 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6888 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.68 1.92 2.255 2.12 ;
        RECT 0.68 0.86 1.39 1.04 ;
        RECT 1.1 0.325 1.39 1.04 ;
        RECT 0.68 1.92 1.01 2.735 ;
        RECT 0.68 0.86 0.85 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.735 -0.085 3.065 1.04 ;
        RECT 0.25 -0.085 0.51 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.805 1.925 3.135 3.415 ;
        RECT 1.605 2.63 2.275 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.445 1.92 2.635 3.075 ;
      RECT 0.25 2.905 1.435 3.075 ;
      RECT 1.18 2.29 1.435 3.075 ;
      RECT 0.25 1.92 0.51 3.075 ;
      RECT 1.18 2.29 2.635 2.46 ;
      RECT 2.425 1.92 2.635 2.46 ;
  END
END scs130lp_a32oi_1

MACRO scs130lp_a32oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32oi_2 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.435 1.425 2.765 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.515 1.425 4.655 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.755 1.195 6.155 1.525 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.895 1.425 2.265 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.275 1.06 1.525 ;
        RECT 0.085 1.21 0.485 1.525 ;
        RECT 0.085 1.21 0.435 1.76 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.92 3.335 2.12 ;
        RECT 3.005 0.605 3.335 2.12 ;
        RECT 1.465 1.075 3.335 1.245 ;
        RECT 1.465 1.92 1.795 2.735 ;
        RECT 1.465 0.605 1.795 1.245 ;
        RECT 1.465 1.695 1.725 2.735 ;
        RECT 0.605 1.695 1.725 1.865 ;
        RECT 0.605 1.695 0.935 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.755 -0.085 6.085 1.025 ;
        RECT 4.895 -0.085 5.225 0.905 ;
        RECT 0.605 -0.085 0.935 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.175 2.095 5.505 3.415 ;
        RECT 3.945 2.26 4.645 3.415 ;
        RECT 2.56 2.63 3.335 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.675 1.755 5.935 3.075 ;
      RECT 4.815 1.92 5.005 3.075 ;
      RECT 3.505 2.29 3.775 3.075 ;
      RECT 3.515 1.92 3.775 3.075 ;
      RECT 0.175 2.905 2.345 3.075 ;
      RECT 2.015 2.29 2.345 3.075 ;
      RECT 1.105 2.035 1.295 3.075 ;
      RECT 0.175 1.93 0.435 3.075 ;
      RECT 2.015 2.29 3.775 2.46 ;
      RECT 3.515 1.92 5.005 2.09 ;
      RECT 4.825 1.755 5.935 1.925 ;
      RECT 3.865 1.075 5.585 1.245 ;
      RECT 5.395 0.255 5.585 1.245 ;
      RECT 3.865 0.605 4.195 1.245 ;
      RECT 3.505 0.265 3.695 1.205 ;
      RECT 4.365 0.265 4.695 0.905 ;
      RECT 2.505 0.265 2.835 0.905 ;
      RECT 2.505 0.265 4.695 0.435 ;
      RECT 0.175 0.87 1.295 1.04 ;
      RECT 1.105 0.265 1.295 1.04 ;
      RECT 1.965 0.265 2.295 0.905 ;
      RECT 0.175 0.315 0.435 1.04 ;
      RECT 1.105 0.265 2.295 0.435 ;
  END
END scs130lp_a32oi_2

MACRO scs130lp_a32oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32oi_4 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.995 1.21 5.715 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.265 1.21 8.005 1.435 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.315 1.21 10.455 1.435 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 3.815 1.435 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 1.845 1.435 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 1.605 6.095 1.875 ;
        RECT 5.885 0.765 6.095 1.875 ;
        RECT 2.25 0.765 6.095 1.04 ;
        RECT 3.18 1.605 3.51 2.735 ;
        RECT 2.32 1.605 2.65 2.735 ;
        RECT 1.46 1.605 1.79 2.735 ;
        RECT 0.6 1.605 0.93 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.84 -0.085 10.17 1.04 ;
        RECT 8.98 -0.085 9.31 0.595 ;
        RECT 8.12 -0.085 8.45 0.595 ;
        RECT 1.39 -0.085 1.72 0.7 ;
        RECT 0.53 -0.085 0.86 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.15 1.945 9.48 3.415 ;
        RECT 8.29 1.945 8.62 3.415 ;
        RECT 7.43 1.945 7.76 3.415 ;
        RECT 6.21 2.395 6.9 3.415 ;
        RECT 5.01 2.445 5.68 3.415 ;
        RECT 4.15 2.395 4.48 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.65 1.605 9.91 3.075 ;
      RECT 8.79 1.605 8.98 3.075 ;
      RECT 7.93 1.605 8.12 3.075 ;
      RECT 7.07 1.605 7.26 3.075 ;
      RECT 5.85 2.045 6.04 3.075 ;
      RECT 4.65 2.045 4.84 3.075 ;
      RECT 0.17 2.905 3.98 3.075 ;
      RECT 3.68 2.045 3.98 3.075 ;
      RECT 2.82 2.045 3.01 3.075 ;
      RECT 1.96 2.045 2.15 3.075 ;
      RECT 1.1 2.045 1.29 3.075 ;
      RECT 0.17 1.825 0.43 3.075 ;
      RECT 3.68 2.045 7.26 2.225 ;
      RECT 7 1.605 7.26 2.225 ;
      RECT 7 1.605 9.91 1.775 ;
      RECT 6.31 0.815 9.67 1.04 ;
      RECT 9.48 0.255 9.67 1.04 ;
      RECT 6.31 0.765 8.81 1.04 ;
      RECT 8.62 0.255 8.81 1.04 ;
      RECT 0.1 0.87 2.08 1.04 ;
      RECT 1.89 0.255 2.08 1.04 ;
      RECT 1.03 0.255 1.22 1.04 ;
      RECT 0.1 0.255 0.36 1.04 ;
      RECT 1.89 0.255 3.87 0.595 ;
      RECT 4.16 0.265 7.93 0.595 ;
  END
END scs130lp_a32oi_4

MACRO scs130lp_a32oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32oi_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.575 0.44 1.935 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.145 1.45 2.755 1.78 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.81 3.235 1.14 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 1.11 1.395 1.78 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 1.12 0.855 1.79 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5089 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.76 1.395 0.93 ;
        RECT 1.065 0.265 1.395 0.93 ;
        RECT 0.79 1.97 1.12 2.715 ;
        RECT 0.125 1.97 1.12 2.14 ;
        RECT 0.125 0.76 0.345 2.14 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.69 -0.085 3.02 0.63 ;
        RECT 0.245 -0.085 0.575 0.58 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.99 2.025 3.24 3.415 ;
        RECT 1.85 2.31 2.18 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.38 1.96 2.71 3.065 ;
      RECT 0.26 2.895 1.65 3.065 ;
      RECT 1.32 1.96 1.65 3.065 ;
      RECT 0.26 2.32 0.59 3.065 ;
      RECT 1.32 1.96 2.71 2.13 ;
  END
END scs130lp_a32oi_lp

MACRO scs130lp_a32oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a32oi_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 0.47 1.765 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.47 2.245 2.12 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.84 2.815 2.49 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.84 1.285 2.12 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.49 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2541 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.49 1.345 0.66 ;
        RECT 1.155 0.33 1.345 0.66 ;
        RECT 0.67 2.3 1 2.71 ;
        RECT 0.635 0.49 0.805 2.47 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.47 -0.085 2.8 0.485 ;
        RECT 0.125 -0.085 0.455 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.55 2.67 2.88 3.415 ;
        RECT 1.61 2.67 1.94 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.16 2.89 1.39 3.06 ;
      RECT 1.18 2.32 1.39 3.06 ;
      RECT 0.16 2.67 0.49 3.06 ;
      RECT 2.2 2.32 2.37 2.81 ;
      RECT 1.18 2.32 2.37 2.49 ;
  END
END scs130lp_a32oi_m

MACRO scs130lp_a41o_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41o_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.77 1.84 1.835 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.01 0.385 2.385 1.835 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.785 0.77 3.215 1.825 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 0.77 3.755 1.835 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 1.08 1.365 1.83 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.28 0.57 0.61 ;
        RECT 0.085 2.385 0.39 3.065 ;
        RECT 0.085 0.28 0.335 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.135 -0.085 3.53 0.6 ;
        RECT 0.74 -0.085 0.995 0.57 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.9 2.345 3.19 3.415 ;
        RECT 2.04 2.345 2.305 3.415 ;
        RECT 0.56 2.385 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.36 2.005 3.655 3.025 ;
      RECT 2.475 2.005 2.73 3.025 ;
      RECT 1.615 2.005 1.87 3.025 ;
      RECT 1.615 2.005 3.655 2.175 ;
      RECT 1.15 2.045 1.445 3.025 ;
      RECT 0.505 2.045 1.445 2.215 ;
      RECT 0.505 1.545 0.895 2.215 ;
      RECT 0.725 0.74 0.895 2.215 ;
      RECT 0.725 0.74 1.415 0.91 ;
      RECT 1.165 0.28 1.415 0.91 ;
      RECT 1.165 0.28 1.8 0.6 ;
  END
END scs130lp_a41o_0

MACRO scs130lp_a41o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41o_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.39 2.345 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 0.39 2.85 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.02 0.39 3.685 1.515 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.855 1.185 4.235 1.515 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.21 1.905 1.435 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.255 0.57 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.855 -0.085 4.135 1.015 ;
        RECT 0.75 -0.085 1.555 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.355 2.025 3.685 3.415 ;
        RECT 2.135 2.025 2.805 3.415 ;
        RECT 0.75 1.945 1.02 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.855 1.685 4.135 3.075 ;
      RECT 2.975 1.685 3.185 3.075 ;
      RECT 1.74 1.685 1.965 3.075 ;
      RECT 1.74 1.685 4.135 1.855 ;
      RECT 1.275 1.605 1.57 3.075 ;
      RECT 0.74 1.605 1.57 1.775 ;
      RECT 0.74 0.87 0.945 1.775 ;
      RECT 0.74 0.87 1.905 1.04 ;
      RECT 1.725 0.255 1.905 1.04 ;
  END
END scs130lp_a41o_1

MACRO scs130lp_a41o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41o_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.345 1.345 4.71 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.475 1.345 4.175 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.975 1.345 3.305 1.75 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 1.345 2.805 1.75 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.345 2.305 1.75 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 0.36 0.835 2.975 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 2.295 -0.085 2.625 0.825 ;
        RECT 1.005 -0.085 1.335 1.175 ;
        RECT 0.145 -0.085 0.43 1.255 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.79 2.27 4.12 3.415 ;
        RECT 2.69 2.27 3.02 3.415 ;
        RECT 1.005 1.845 1.335 3.415 ;
        RECT 0.145 1.815 0.43 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.81 1.92 2.08 3.075 ;
      RECT 1.665 0.255 1.835 2.1 ;
      RECT 1.025 1.345 1.835 1.675 ;
      RECT 1.505 0.255 1.835 1.675 ;
      RECT 1.505 0.995 4.55 1.165 ;
      RECT 4.22 0.255 4.55 1.165 ;
      RECT 1.505 0.255 2.08 1.165 ;
      RECT 4.29 1.92 4.55 3.075 ;
      RECT 3.26 1.92 3.59 3.075 ;
      RECT 2.3 1.92 2.52 3.075 ;
      RECT 2.3 1.92 4.55 2.1 ;
  END
END scs130lp_a41o_2

MACRO scs130lp_a41o_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41o_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.89 1.21 4.7 1.585 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.87 1.185 5.17 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.365 1.21 6.085 1.52 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.395 1.21 7.58 1.575 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.765 1.195 3.72 1.535 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.555 1.755 1.78 3.075 ;
        RECT 0.1 1.055 1.78 1.225 ;
        RECT 1.555 0.255 1.78 1.225 ;
        RECT 0.1 1.755 1.78 1.925 ;
        RECT 0.695 1.755 0.885 3.075 ;
        RECT 0.695 0.255 0.885 1.225 ;
        RECT 0.1 1.055 0.42 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.825 -0.085 7.155 0.7 ;
        RECT 2.775 -0.085 3.105 0.515 ;
        RECT 1.95 -0.085 2.21 1.105 ;
        RECT 1.055 -0.085 1.385 0.885 ;
        RECT 0.195 -0.085 0.525 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.35 2.095 6.68 3.415 ;
        RECT 5.49 2.095 5.82 3.415 ;
        RECT 4.605 2.095 4.935 3.415 ;
        RECT 3.725 2.095 4.055 3.415 ;
        RECT 1.95 1.815 2.235 3.415 ;
        RECT 1.055 2.095 1.385 3.415 ;
        RECT 0.195 2.095 0.525 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.535 0.87 7.585 1.04 ;
      RECT 7.325 0.255 7.585 1.04 ;
      RECT 5.535 0.765 6.655 1.04 ;
      RECT 6.405 0.255 6.655 1.04 ;
      RECT 6.85 1.755 7.11 3.075 ;
      RECT 5.99 1.755 6.18 3.075 ;
      RECT 5.11 1.755 5.32 3.075 ;
      RECT 4.225 1.755 4.415 3.075 ;
      RECT 2.435 2.905 3.555 3.075 ;
      RECT 3.365 1.755 3.555 3.075 ;
      RECT 2.435 2.045 2.695 3.075 ;
      RECT 3.365 1.755 7.11 1.925 ;
      RECT 4.155 0.765 5.345 1.015 ;
      RECT 4.155 0.255 4.425 1.015 ;
      RECT 3.295 0.255 4.425 0.505 ;
      RECT 2.865 1.705 3.195 2.735 ;
      RECT 2.405 1.705 3.195 1.875 ;
      RECT 2.405 0.255 2.595 1.875 ;
      RECT 0.59 1.405 2.595 1.575 ;
      RECT 2.38 0.255 2.595 1.575 ;
      RECT 2.38 0.685 3.985 1.015 ;
      RECT 2.38 0.255 2.605 1.015 ;
      RECT 4.595 0.265 6.235 0.595 ;
  END
END scs130lp_a41o_4

MACRO scs130lp_a41o_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41o_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 1.075 2.32 1.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.42 0.44 1.795 1.435 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.615 0.44 1.21 1.435 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.825 0.435 1.495 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.075 2.99 1.745 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.875 0.265 4.205 3.065 ;
        RECT 3.835 0.265 4.205 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.045 -0.085 3.375 0.545 ;
        RECT 0.185 -0.085 0.435 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.345 2.275 3.675 3.415 ;
        RECT 1.705 2.275 2.035 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.785 1.925 3.115 3.065 ;
      RECT 2.785 1.925 3.655 2.095 ;
      RECT 3.325 0.725 3.655 2.095 ;
      RECT 2.255 0.725 3.655 0.895 ;
      RECT 2.255 0.265 2.585 0.895 ;
      RECT 2.255 1.925 2.585 3.065 ;
      RECT 1.175 1.675 1.505 3.065 ;
      RECT 0.115 1.675 0.445 3.065 ;
      RECT 1.175 1.925 2.585 2.095 ;
      RECT 0.115 1.675 1.505 1.845 ;
  END
END scs130lp_a41o_lp

MACRO scs130lp_a41o_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41o_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.47 1.775 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.47 2.315 2.12 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.84 2.855 2.12 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.345 0.84 3.685 2.12 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 1.21 1.285 2.215 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.265 0.575 0.595 ;
        RECT 0.155 0.265 0.345 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.09 -0.085 3.42 0.485 ;
        RECT 0.795 -0.085 1.005 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.825 2.65 3.035 3.415 ;
        RECT 1.905 2.71 2.235 3.415 ;
        RECT 0.525 2.845 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.255 2.3 3.465 2.85 ;
      RECT 2.415 2.3 2.605 2.85 ;
      RECT 1.535 2.3 1.725 2.85 ;
      RECT 1.535 2.3 3.465 2.47 ;
      RECT 1.105 2.395 1.315 2.85 ;
      RECT 0.525 2.395 1.315 2.565 ;
      RECT 0.525 0.775 0.695 2.565 ;
      RECT 0.525 0.775 1.415 0.945 ;
      RECT 1.225 0.345 1.415 0.945 ;
  END
END scs130lp_a41o_m

MACRO scs130lp_a41oi_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41oi_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.99 0.825 1.36 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 0.825 1.855 1.84 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 0.825 2.355 1.84 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.995 3.275 1.84 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.825 0.45 1.495 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3208 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.62 0.28 2.415 0.655 ;
        RECT 0.62 0.28 0.82 1.855 ;
        RECT 0.425 1.685 0.72 3.055 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.715 -0.085 3.045 0.61 ;
        RECT 0.245 -0.085 0.45 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.175 2.375 2.445 3.415 ;
        RECT 1.32 2.375 1.575 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.615 2.025 2.905 3.055 ;
      RECT 1.745 2.025 2.005 3.055 ;
      RECT 0.89 2.025 1.15 3.055 ;
      RECT 0.89 2.025 2.905 2.205 ;
  END
END scs130lp_a41oi_0

MACRO scs130lp_a41oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41oi_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.92 1.185 3.275 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.27 1.175 2.75 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.175 2.06 1.75 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.04 1.175 1.355 1.75 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.185 0.405 1.515 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7791 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.185 0.835 3.265 1.005 ;
        RECT 2.935 0.265 3.265 1.005 ;
        RECT 0.185 1.695 0.87 1.865 ;
        RECT 0.575 0.835 0.87 1.865 ;
        RECT 0.185 0.835 0.87 1.015 ;
        RECT 0.185 1.695 0.445 3.075 ;
        RECT 0.185 0.265 0.445 1.015 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 0.615 -0.085 1.395 0.665 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.485 2.26 2.815 3.415 ;
        RECT 1.075 2.375 1.935 3.415 ;
        RECT 1.455 2.265 1.935 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.985 1.92 3.265 3.075 ;
      RECT 2.105 1.92 2.315 3.075 ;
      RECT 0.615 2.035 0.905 3.075 ;
      RECT 0.615 2.035 1.285 2.205 ;
      RECT 0.615 2.035 2.315 2.095 ;
      RECT 1.635 1.92 3.265 2.09 ;
      RECT 1.115 1.925 3.265 2.09 ;
  END
END scs130lp_a41oi_1

MACRO scs130lp_a41oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41oi_2 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.21 1.9 1.61 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.97 1.425 3.685 1.83 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.105 1.375 4.785 1.545 ;
        RECT 4.4 1.21 4.73 1.545 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.25 1.425 6.155 1.75 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.805 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8232 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.07 1.425 2.8 1.95 ;
        RECT 2.07 0.595 2.33 1.95 ;
        RECT 0.975 1.78 2.8 1.95 ;
        RECT 0.67 0.87 2.33 1.04 ;
        RECT 2 0.595 2.33 1.04 ;
        RECT 0.905 1.89 1.235 2.725 ;
        RECT 0.67 0.255 0.86 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.26 -0.085 5.59 0.915 ;
        RECT 1.03 -0.085 1.36 0.7 ;
        RECT 0.17 -0.085 0.5 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.26 2.265 5.59 3.415 ;
        RECT 4.315 2.055 4.645 3.415 ;
        RECT 2.86 2.505 3.7 3.415 ;
        RECT 1.845 2.46 2.175 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.91 1.085 6.02 1.255 ;
      RECT 5.76 0.325 6.02 1.255 ;
      RECT 3.9 0.595 4.23 1.205 ;
      RECT 4.91 0.325 5.09 1.255 ;
      RECT 3.9 0.87 5.09 1.04 ;
      RECT 4.9 0.325 5.09 1.04 ;
      RECT 5.76 1.925 6.02 3.075 ;
      RECT 4.83 1.925 5.09 3.075 ;
      RECT 3.87 1.715 4.13 3.075 ;
      RECT 2.36 2.12 2.69 3.075 ;
      RECT 0.475 2.895 1.665 3.075 ;
      RECT 1.405 2.12 1.665 3.075 ;
      RECT 1.335 2.885 1.665 3.075 ;
      RECT 0.475 1.92 0.735 3.075 ;
      RECT 2.36 2.12 4.13 2.325 ;
      RECT 3.855 1.715 4.13 2.325 ;
      RECT 1.405 2.12 4.13 2.29 ;
      RECT 4.83 1.925 6.02 2.095 ;
      RECT 4.83 1.715 5.08 3.075 ;
      RECT 3.855 1.715 5.08 1.885 ;
      RECT 2.86 0.255 3.19 0.915 ;
      RECT 4.4 0.255 4.73 0.7 ;
      RECT 2.86 0.255 4.73 0.425 ;
      RECT 2.5 1.085 3.69 1.255 ;
      RECT 3.36 0.595 3.69 1.255 ;
      RECT 2.5 0.255 2.69 1.255 ;
      RECT 1.55 0.255 1.83 0.7 ;
      RECT 1.55 0.255 2.69 0.425 ;
  END
END scs130lp_a41oi_2

MACRO scs130lp_a41oi_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41oi_4 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.405 4.095 1.575 ;
        RECT 2.555 1.21 3.205 1.575 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.625 1.195 5.975 1.585 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.185 1.355 8.215 1.585 ;
        RECT 6.185 1.315 7.535 1.585 ;
        RECT 7.345 1.155 7.535 1.585 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.425 1.2 10.455 1.585 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.21 1.825 1.435 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.4 1.745 4.455 1.935 ;
        RECT 4.265 1.065 4.455 1.935 ;
        RECT 3.64 1.065 4.455 1.235 ;
        RECT 3.64 0.595 3.97 1.235 ;
        RECT 0.595 0.855 3.97 1.04 ;
        RECT 1.455 0.815 3.97 1.04 ;
        RECT 0.54 1.605 1.815 1.79 ;
        RECT 1.4 1.605 1.73 2.735 ;
        RECT 1.455 0.255 1.645 1.04 ;
        RECT 0.54 1.605 0.87 2.735 ;
        RECT 0.595 0.255 0.785 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.425 -0.085 9.755 0.69 ;
        RECT 8.565 -0.085 8.895 0.69 ;
        RECT 1.815 -0.085 2.145 0.645 ;
        RECT 0.955 -0.085 1.285 0.685 ;
        RECT 0.095 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.41 2.105 9.74 3.415 ;
        RECT 8.55 2.105 8.88 3.415 ;
        RECT 7.17 2.105 8.02 3.415 ;
        RECT 6.31 2.105 6.64 3.415 ;
        RECT 5.37 2.105 5.7 3.415 ;
        RECT 4.5 2.455 4.72 3.415 ;
        RECT 3.16 2.465 3.83 3.415 ;
        RECT 2.28 2.455 2.61 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.215 0.86 10.185 1.03 ;
      RECT 9.925 0.315 10.185 1.03 ;
      RECT 9.065 0.315 9.255 1.03 ;
      RECT 8.215 0.255 8.395 1.03 ;
      RECT 7.345 0.255 7.535 0.645 ;
      RECT 6.475 0.255 6.675 0.645 ;
      RECT 6.475 0.255 8.395 0.425 ;
      RECT 9.91 1.755 10.17 3.075 ;
      RECT 9.05 1.755 9.24 3.075 ;
      RECT 8.19 1.755 8.38 3.075 ;
      RECT 6.81 1.755 7 3.075 ;
      RECT 5.88 1.755 6.14 3.075 ;
      RECT 4.89 1.755 5.13 3.075 ;
      RECT 4 2.105 4.33 3.075 ;
      RECT 2.78 2.105 2.99 3.075 ;
      RECT 0.11 2.905 2.11 3.075 ;
      RECT 1.9 2.105 2.11 3.075 ;
      RECT 1.04 1.96 1.23 3.075 ;
      RECT 0.11 1.825 0.37 3.075 ;
      RECT 1.9 2.105 5.13 2.285 ;
      RECT 4.86 1.755 5.13 2.285 ;
      RECT 4.86 1.755 10.17 1.925 ;
      RECT 7.705 0.615 8.035 1.145 ;
      RECT 6.845 0.615 7.175 1.145 ;
      RECT 4.65 0.815 7.175 1.025 ;
      RECT 4.65 0.815 8.035 0.985 ;
      RECT 4.65 0.595 4.9 1.025 ;
      RECT 4.15 0.255 4.48 0.895 ;
      RECT 5.07 0.255 6.14 0.645 ;
      RECT 2.35 0.255 3.47 0.645 ;
      RECT 2.35 0.255 6.14 0.425 ;
  END
END scs130lp_a41oi_4

MACRO scs130lp_a41oi_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41oi_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 1.12 2.32 1.79 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.45 0.44 1.795 1.79 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.45 1.24 1.78 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.81 0.835 1.14 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.12 2.89 1.79 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.785 2.025 3.24 3.065 ;
        RECT 3.07 0.77 3.24 3.065 ;
        RECT 2.045 0.77 3.24 0.94 ;
        RECT 2.045 0.265 2.445 0.94 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.905 -0.085 3.235 0.59 ;
        RECT 0.395 -0.085 0.725 0.63 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.705 2.32 2.035 3.415 ;
        RECT 0.645 2.32 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.255 1.97 2.585 3.065 ;
      RECT 1.175 1.97 1.505 3.065 ;
      RECT 0.115 1.97 0.445 3.065 ;
      RECT 0.115 1.97 2.585 2.14 ;
  END
END scs130lp_a41oi_lp

MACRO scs130lp_a41oi_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_a41oi_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.21 1.325 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.47 1.89 2.12 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.435 0.84 2.725 2.185 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 0.84 3.205 2.49 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.615 1.21 0.805 2.86 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3507 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 1.315 1.01 ;
        RECT 1.105 0.345 1.315 1.01 ;
        RECT 0.155 0.84 0.435 2.965 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.665 -0.085 2.995 0.485 ;
        RECT 0.675 -0.085 0.885 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.255 2.785 2.445 3.415 ;
        RECT 1.395 2.785 1.605 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.825 2.435 2.035 2.965 ;
      RECT 0.985 2.435 1.175 2.945 ;
      RECT 2.625 2.695 2.955 2.905 ;
      RECT 2.625 2.435 2.795 2.905 ;
      RECT 0.985 2.435 2.795 2.605 ;
  END
END scs130lp_a41oi_m

MACRO scs130lp_and2_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2_0 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.185 0.545 2.23 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.075 1.535 1.395 2.205 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.935 2.385 2.315 3.055 ;
        RECT 2.065 0.28 2.315 3.055 ;
        RECT 1.52 0.28 2.315 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.065 -0.085 1.35 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.15 2.385 1.765 3.415 ;
        RECT 0.275 2.44 0.545 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.715 2.44 0.98 2.77 ;
      RECT 0.715 0.845 0.895 2.77 ;
      RECT 1.565 0.845 1.895 1.435 ;
      RECT 0.3 0.845 1.895 1.015 ;
      RECT 0.3 0.28 0.605 1.015 ;
  END
END scs130lp_and2_0

MACRO scs130lp_and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.49 0.865 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.49 1.435 1.75 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5817 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 0.255 2.315 3.075 ;
        RECT 1.75 0.255 2.315 0.98 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.21 -0.085 1.58 0.98 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.545 2.26 1.875 3.415 ;
        RECT 0.42 1.955 0.75 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.92 1.92 1.25 2.285 ;
      RECT 0.92 1.92 1.875 2.09 ;
      RECT 1.625 1.15 1.875 2.09 ;
      RECT 0.42 1.15 1.875 1.32 ;
      RECT 0.42 0.7 0.75 1.32 ;
  END
END scs130lp_and2_1

MACRO scs130lp_and2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2_2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.035 0.435 1.86 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.125 1.005 1.43 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.94 1.815 3.075 ;
        RECT 1.635 0.255 1.815 3.075 ;
        RECT 1.575 0.255 1.815 1.09 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.985 -0.085 2.265 1.09 ;
        RECT 1.03 -0.085 1.36 0.525 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.985 1.815 2.265 3.415 ;
        RECT 1.015 1.945 1.36 3.415 ;
        RECT 0.12 2.03 0.45 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.62 1.6 0.845 2.36 ;
      RECT 0.62 1.6 1.465 1.77 ;
      RECT 1.235 1.27 1.465 1.77 ;
      RECT 1.235 0.695 1.405 1.77 ;
      RECT 0.19 0.695 1.405 0.865 ;
      RECT 0.19 0.28 0.52 0.865 ;
  END
END scs130lp_and2_2

MACRO scs130lp_and2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2_4 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.325 0.455 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.325 1.02 1.75 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.775 3.26 1.945 ;
        RECT 2.855 1.065 3.26 1.945 ;
        RECT 1.53 1.065 3.26 1.235 ;
        RECT 2.39 1.775 2.58 3.075 ;
        RECT 2.39 0.255 2.58 1.235 ;
        RECT 1.53 1.775 1.72 3.075 ;
        RECT 1.53 0.255 1.72 1.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.75 -0.085 3.08 0.885 ;
        RECT 1.89 -0.085 2.22 0.885 ;
        RECT 0.955 -0.085 1.285 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.75 2.115 3.08 3.415 ;
        RECT 1.89 2.115 2.22 3.415 ;
        RECT 0.99 2.27 1.32 3.415 ;
        RECT 0.095 1.92 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.595 1.93 0.785 3.075 ;
      RECT 0.595 1.93 1.36 2.1 ;
      RECT 1.19 0.985 1.36 2.1 ;
      RECT 1.19 1.405 2.685 1.605 ;
      RECT 0.095 0.985 1.36 1.155 ;
      RECT 0.095 0.255 0.425 1.155 ;
  END
END scs130lp_and2_4

MACRO scs130lp_and2_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 0.35 1.845 0.68 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.48 1.315 2.15 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.44 3.235 2.89 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.015 -0.085 2.345 0.9 ;
        RECT 0.43 -0.085 0.76 1.31 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.83 2.32 2.16 3.415 ;
        RECT 0.25 2.32 0.58 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.04 2.32 1.655 2.78 ;
      RECT 1.485 0.85 1.655 2.78 ;
      RECT 2.025 1.07 2.355 1.74 ;
      RECT 1.25 1.14 2.355 1.31 ;
      RECT 1.25 0.85 1.655 1.31 ;
  END
END scs130lp_and2_lp

MACRO scs130lp_and2_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2_lp2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.85 1.165 2.275 1.835 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.165 1.435 1.495 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 2.025 0.61 3.065 ;
        RECT 0.125 0.265 0.52 0.635 ;
        RECT 0.125 0.265 0.355 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.98 -0.085 1.31 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.9 2.025 2.23 3.415 ;
        RECT 0.81 2.025 1.14 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.34 1.675 1.67 3.065 ;
      RECT 0.535 1.675 1.67 1.845 ;
      RECT 0.535 0.815 0.865 1.845 ;
      RECT 0.535 0.815 2.13 0.985 ;
      RECT 1.8 0.265 2.13 0.985 ;
  END
END scs130lp_and2_lp2

MACRO scs130lp_and2_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.435 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.265 1.045 0.64 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.575 0.47 1.765 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.125 0.82 1.395 1.15 ;
        RECT 1.225 -0.085 1.395 1.15 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.125 2.095 1.335 3.415 ;
        RECT 0.17 2.095 0.38 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.615 0.82 0.945 3.025 ;
      RECT 0.13 0.82 0.945 1.03 ;
  END
END scs130lp_and2_m

MACRO scs130lp_and2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2b_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 0.765 0.875 1.095 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 2.32 1.845 3.075 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.455 1.695 2.795 3.075 ;
        RECT 2.49 0.255 2.795 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.835 -0.085 2.32 1.015 ;
        RECT 0.555 -0.085 0.855 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.015 1.765 2.285 3.415 ;
        RECT 1.865 1.765 2.285 2.15 ;
        RECT 0.71 1.87 1.095 2.15 ;
        RECT 0.71 1.87 0.885 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.395 1.185 1.695 2.15 ;
      RECT 1.395 1.185 2.32 1.515 ;
      RECT 1.395 0.695 1.575 2.15 ;
      RECT 1.045 0.695 1.575 1.025 ;
      RECT 0.095 1.335 0.54 2.21 ;
      RECT 0.095 1.335 1.225 1.665 ;
      RECT 0.095 0.28 0.385 2.21 ;
  END
END scs130lp_and2b_1

MACRO scs130lp_and2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2b_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.185 0.92 1.75 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 1.2 2.735 1.455 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.09 0.875 1.56 1.125 ;
        RECT 1.09 0.875 1.315 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.74 -0.085 2.07 0.365 ;
        RECT 0.72 -0.085 1.05 0.365 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.61 1.965 2.94 3.415 ;
        RECT 1.485 1.965 2.08 3.415 ;
        RECT 0.6 1.92 0.92 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.25 1.625 2.44 2.21 ;
      RECT 1.485 1.625 3.16 1.795 ;
      RECT 2.905 0.725 3.16 1.795 ;
      RECT 1.485 1.345 1.735 1.795 ;
      RECT 2.61 0.725 3.16 1.03 ;
      RECT 0.09 1.92 0.43 2.21 ;
      RECT 0.09 0.535 0.26 2.21 ;
      RECT 0.09 0.535 0.52 1.015 ;
      RECT 0.09 0.535 2.43 0.705 ;
      RECT 2.26 0.255 2.815 0.555 ;
  END
END scs130lp_and2b_2

MACRO scs130lp_and2b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2b_4 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.19 0.88 2.205 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.83 1.345 3.215 1.76 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.05 1.075 2.31 1.245 ;
        RECT 2.12 0.255 2.31 1.245 ;
        RECT 1.05 1.815 2.3 2.145 ;
        RECT 1.23 0.255 1.45 1.245 ;
        RECT 1.05 1.075 1.285 2.145 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.55 -0.085 2.88 0.815 ;
        RECT 1.62 -0.085 1.95 0.895 ;
        RECT 0.76 -0.085 1.06 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.415 2.78 3.745 3.415 ;
        RECT 2.515 2.78 2.845 3.415 ;
        RECT 1.62 2.78 1.95 3.415 ;
        RECT 0.76 2.78 1.09 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.48 1.93 3.255 2.26 ;
      RECT 2.48 0.995 2.66 2.26 ;
      RECT 1.495 1.415 2.66 1.645 ;
      RECT 2.48 0.995 3.745 1.165 ;
      RECT 3.415 0.255 3.745 1.165 ;
      RECT 0.175 2.43 3.715 2.61 ;
      RECT 3.545 1.375 3.715 2.61 ;
      RECT 0.175 0.72 0.425 2.61 ;
      RECT 3.385 1.375 3.715 1.545 ;
      RECT 0.175 0.72 0.565 1.02 ;
  END
END scs130lp_and2b_4

MACRO scs130lp_and2b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2b_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.035 2.855 1.41 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.32 1.605 1.795 2.15 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.44 0.57 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.095 -0.085 2.425 0.675 ;
        RECT 1.055 -0.085 1.385 1.075 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.115 2.115 2.445 3.415 ;
        RECT 0.85 2.68 1.18 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.77 1.605 3.1 3.065 ;
      RECT 1.975 1.605 3.245 1.935 ;
      RECT 3.075 0.295 3.245 1.935 ;
      RECT 2.915 0.295 3.245 0.675 ;
      RECT 1.585 2.33 1.915 3.065 ;
      RECT 0.75 2.33 1.915 2.5 ;
      RECT 0.75 1.255 1.08 2.5 ;
      RECT 0.75 1.255 2.345 1.425 ;
      RECT 2.015 0.905 2.345 1.425 ;
  END
END scs130lp_and2b_lp

MACRO scs130lp_and2b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and2b_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.52 0.84 1.285 1.38 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.87 0.84 2.245 1.825 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 0.345 2.725 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.085 -0.085 2.275 0.545 ;
        RECT 0.565 -0.085 0.895 0.6 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.005 2.155 2.335 3.415 ;
        RECT 0.855 2.095 1.065 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.495 2.855 1.825 3.025 ;
      RECT 1.495 2.155 1.69 3.025 ;
      RECT 1.52 0.405 1.69 3.025 ;
      RECT 1.315 2.155 1.69 2.365 ;
      RECT 1.235 0.405 1.69 0.615 ;
      RECT 0.17 2.025 0.675 2.235 ;
      RECT 0.17 0.33 0.34 2.235 ;
      RECT 0.17 1.575 1.34 1.745 ;
      RECT 0.17 0.33 0.385 0.66 ;
  END
END scs130lp_and2b_m

MACRO scs130lp_and3_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.495 0.84 0.86 1.835 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 1.17 1.36 1.915 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.17 1.895 2.18 ;
        RECT 1.53 1.17 1.895 1.925 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2873 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.43 2.395 2.795 3.065 ;
        RECT 2.525 0.345 2.795 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.48 -0.085 2.355 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.655 2.395 2.26 3.415 ;
        RECT 0.795 2.46 1.055 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.225 2.46 1.485 2.79 ;
      RECT 0.155 2.095 0.625 2.79 ;
      RECT 1.225 2.095 1.415 2.79 ;
      RECT 0.155 2.095 1.415 2.265 ;
      RECT 0.155 0.37 0.325 2.79 ;
      RECT 2.105 0.83 2.355 1.625 ;
      RECT 1.09 0.83 2.355 1 ;
      RECT 1.09 0.37 1.26 1 ;
      RECT 0.155 0.37 1.26 0.67 ;
  END
END scs130lp_and3_0

MACRO scs130lp_and3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.485 1.105 0.815 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.105 1.34 1.435 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 2.355 1.775 2.94 ;
        RECT 1.595 1.105 1.775 2.94 ;
        RECT 1.575 1.105 1.775 1.52 ;
        RECT 1.51 1.105 1.775 1.455 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.495 0.255 2.795 3.075 ;
        RECT 2.295 0.255 2.795 1.125 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.74 -0.085 2.07 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.945 1.81 2.325 3.415 ;
        RECT 0.735 1.945 1.015 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.185 1.605 1.425 2.21 ;
      RECT 0.145 1.605 0.565 2.21 ;
      RECT 0.145 1.605 1.425 1.775 ;
      RECT 1.945 1.305 2.325 1.635 ;
      RECT 0.145 0.31 0.315 2.21 ;
      RECT 1.945 0.765 2.125 1.635 ;
      RECT 0.145 0.765 2.125 0.935 ;
      RECT 0.145 0.31 0.62 0.935 ;
  END
END scs130lp_and3_1

MACRO scs130lp_and3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3_2 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.11 1.015 0.44 1.525 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.125 0.9 1.455 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.185 1.44 1.515 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.815 2.33 3.075 ;
        RECT 2.15 0.255 2.33 3.075 ;
        RECT 2.065 0.255 2.33 1.095 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.5 -0.085 2.76 1.085 ;
        RECT 1.445 -0.085 1.775 0.505 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.5 1.815 2.76 3.415 ;
        RECT 1.46 2.045 1.855 3.415 ;
        RECT 0.56 2.045 0.82 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.99 1.705 1.29 2.3 ;
      RECT 0.095 1.705 0.39 2.3 ;
      RECT 0.095 1.705 1.865 1.875 ;
      RECT 1.695 0.675 1.865 1.875 ;
      RECT 1.695 1.275 1.98 1.605 ;
      RECT 0.165 0.675 1.865 0.845 ;
      RECT 0.165 0.255 0.495 0.845 ;
  END
END scs130lp_and3_2

MACRO scs130lp_and3_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3_4 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.21 0.805 1.515 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 1.21 1.34 1.54 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.81 1.54 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.32 1.755 4.225 1.925 ;
        RECT 3.995 0.39 4.225 1.925 ;
        RECT 2.32 1.065 4.225 1.235 ;
        RECT 3.18 1.755 3.37 3.075 ;
        RECT 3.18 0.255 3.37 1.235 ;
        RECT 2.32 1.755 2.51 3.075 ;
        RECT 2.32 0.255 2.51 1.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.54 -0.085 3.825 0.895 ;
        RECT 2.68 -0.085 3.01 0.895 ;
        RECT 1.745 -0.085 2.075 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.54 2.095 3.87 3.415 ;
        RECT 2.68 2.095 3.01 3.415 ;
        RECT 1.765 2.05 2.095 3.415 ;
        RECT 0.815 2.105 1.145 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.35 1.71 1.595 3.075 ;
      RECT 0.345 1.71 0.615 3.075 ;
      RECT 0.345 1.71 1.595 1.925 ;
      RECT 0.345 1.71 2.15 1.88 ;
      RECT 1.98 0.87 2.15 1.88 ;
      RECT 1.98 1.415 3.815 1.585 ;
      RECT 0.345 0.87 2.15 1.04 ;
      RECT 0.345 0.255 0.675 1.04 ;
  END
END scs130lp_and3_4

MACRO scs130lp_and3_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3_lp 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.855 0.435 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.965 1.2 1.315 1.87 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.2 1.865 1.87 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.33 2.06 2.785 3.065 ;
        RECT 2.615 0.265 2.785 3.065 ;
        RECT 2.045 0.265 2.785 0.67 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.535 -0.085 1.865 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.76 2.06 2.09 3.415 ;
        RECT 0.7 2.4 1.03 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.23 2.05 1.56 3.065 ;
      RECT 0.17 2.05 0.5 3.065 ;
      RECT 0.17 2.05 1.56 2.22 ;
      RECT 0.615 0.265 0.785 2.22 ;
      RECT 2.105 0.85 2.435 1.52 ;
      RECT 0.615 0.85 2.435 1.02 ;
      RECT 0.325 0.265 0.785 0.675 ;
  END
END scs130lp_and3_lp

MACRO scs130lp_and3_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.43 1.51 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.96 0.47 1.285 1.435 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 0.84 1.765 1.75 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 0.345 2.245 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.605 -0.085 1.815 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.645 2.065 1.815 3.415 ;
        RECT 1.565 2.065 1.815 2.395 ;
        RECT 0.725 2.065 0.915 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.135 2.825 1.465 2.995 ;
      RECT 1.135 1.935 1.345 2.995 ;
      RECT 0.215 1.715 0.545 2.205 ;
      RECT 1.135 1.715 1.305 2.995 ;
      RECT 0.215 1.715 1.305 1.885 ;
      RECT 0.61 0.33 0.78 1.885 ;
      RECT 0.275 0.33 0.78 0.66 ;
  END
END scs130lp_and3_m

MACRO scs130lp_and3b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3b_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.81 0.395 2.215 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.385 1.86 1.485 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 0.385 2.34 1.435 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.88 1.85 3.275 3.075 ;
        RECT 3.06 0.255 3.275 3.075 ;
        RECT 2.99 0.255 3.275 1.095 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.51 -0.085 2.82 1.095 ;
        RECT 0.095 -0.085 0.395 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.295 2.015 2.66 3.415 ;
        RECT 1.355 2.015 1.685 3.415 ;
        RECT 0.095 2.605 0.395 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.855 1.675 2.125 2.21 ;
      RECT 0.925 1.675 1.185 2.21 ;
      RECT 0.925 1.675 2.7 1.845 ;
      RECT 2.53 1.34 2.7 1.845 ;
      RECT 1.22 0.28 1.395 1.845 ;
      RECT 2.53 1.34 2.89 1.67 ;
      RECT 1.065 0.28 1.395 0.585 ;
      RECT 0.565 2.605 0.855 2.935 ;
      RECT 0.565 0.28 0.755 2.935 ;
      RECT 0.565 0.765 1.05 1.435 ;
      RECT 0.565 0.28 0.855 1.435 ;
  END
END scs130lp_and3b_1

MACRO scs130lp_and3b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3b_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.505 1.21 0.92 1.76 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.535 1.13 3.23 1.485 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 1.13 2.365 1.545 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.885 1.475 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.69 -0.085 2.02 0.375 ;
        RECT 0.62 -0.085 0.95 0.375 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.895 1.995 3.225 3.415 ;
        RECT 1.645 2.095 1.925 3.415 ;
        RECT 0.655 1.93 0.945 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.41 0.73 3.67 2.2 ;
      RECT 2.405 1.715 2.715 2.2 ;
      RECT 1.645 1.715 2.715 1.925 ;
      RECT 3.4 0.73 3.67 1.825 ;
      RECT 2.545 1.655 3.67 1.825 ;
      RECT 1.645 1.295 1.855 1.925 ;
      RECT 0.095 1.93 0.485 2.2 ;
      RECT 0.095 0.545 0.325 2.2 ;
      RECT 0.095 0.545 0.425 1.04 ;
      RECT 1.645 0.545 3.23 0.87 ;
      RECT 0.095 0.545 3.23 0.715 ;
      RECT 3.045 0.255 3.375 0.56 ;
  END
END scs130lp_and3b_2

MACRO scs130lp_and3b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3b_4 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.47 0.805 2.12 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.425 1.345 3.695 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.965 1.345 3.255 1.75 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.075 2.455 1.245 ;
        RECT 2.265 0.255 2.455 1.245 ;
        RECT 0.985 1.815 2.445 2.145 ;
        RECT 1.365 0.255 1.595 1.245 ;
        RECT 0.985 1.075 1.155 2.145 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 2.695 -0.085 3.025 0.825 ;
        RECT 1.765 -0.085 2.095 0.895 ;
        RECT 0.975 -0.085 1.195 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.56 2.78 3.89 3.415 ;
        RECT 2.625 2.78 2.955 3.415 ;
        RECT 1.765 2.655 2.095 3.415 ;
        RECT 0.905 2.655 1.235 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.205 1.815 4.69 3.075 ;
      RECT 4.52 0.255 4.69 3.075 ;
      RECT 2.625 1.93 3.4 2.26 ;
      RECT 2.625 0.995 2.795 2.26 ;
      RECT 1.335 1.425 2.795 1.595 ;
      RECT 2.625 0.995 4.69 1.165 ;
      RECT 3.33 0.255 4.69 1.165 ;
      RECT 2.265 2.43 4.035 2.61 ;
      RECT 3.865 1.335 4.035 2.61 ;
      RECT 0.205 2.315 2.455 2.485 ;
      RECT 0.205 0.7 0.455 2.485 ;
      RECT 3.865 1.335 4.34 1.645 ;
  END
END scs130lp_and3b_4

MACRO scs130lp_and3b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3b_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.905 0.455 1.78 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.17 2.345 1.84 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.17 2.915 1.84 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.445 2.025 4.195 3.065 ;
        RECT 3.665 1.18 4.195 3.065 ;
        RECT 3.665 0.265 3.995 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 2.71 -0.085 3.04 0.64 ;
        RECT 0.115 -0.085 0.445 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.81 2.37 3.14 3.415 ;
        RECT 1.75 2.37 2.08 3.415 ;
        RECT 0.13 2.02 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.28 2.02 2.61 3.065 ;
      RECT 1.22 2.02 1.55 3.065 ;
      RECT 1.22 2.02 3.265 2.19 ;
      RECT 3.095 0.82 3.265 2.19 ;
      RECT 3.095 0.82 3.485 1.49 ;
      RECT 1.5 0.82 3.485 0.99 ;
      RECT 1.5 0.265 1.83 0.99 ;
      RECT 0.66 2.02 0.99 3.06 ;
      RECT 0.82 0.265 0.99 3.06 ;
      RECT 0.82 1.17 1.385 1.84 ;
      RECT 0.82 0.265 1.265 1.84 ;
  END
END scs130lp_and3b_lp

MACRO scs130lp_and3b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and3b_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.49 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.47 1.98 1.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.35 0.84 2.725 1.855 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 0.375 3.265 2.49 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.395 -0.085 2.725 0.515 ;
        RECT 0.155 -0.085 0.365 0.575 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.49 2.125 2.7 3.415 ;
        RECT 1.57 2.125 1.76 3.415 ;
        RECT 0.155 2.67 0.345 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.98 2.855 2.31 3.025 ;
      RECT 1.98 1.775 2.17 3.025 ;
      RECT 1.12 1.945 1.39 2.325 ;
      RECT 1.22 0.405 1.39 2.325 ;
      RECT 1.22 1.775 2.17 1.945 ;
      RECT 1.06 0.405 1.39 0.615 ;
      RECT 0.585 0.33 0.795 3 ;
      RECT 0.585 0.795 1.04 1.465 ;
  END
END scs130lp_and3b_m

MACRO scs130lp_and4_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.83 0.435 2.215 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.945 1.16 1.335 1.88 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.505 1.17 1.825 1.84 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 1.16 2.325 2.21 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.84 2.37 3.275 3.04 ;
        RECT 2.985 0.32 3.275 3.04 ;
        RECT 2.695 0.32 3.275 0.65 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.89 -0.085 2.525 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.995 2.38 2.67 3.415 ;
        RECT 1.085 2.435 1.385 3.415 ;
        RECT 0.19 2.435 0.485 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.655 2.06 0.915 2.765 ;
      RECT 1.555 2.06 1.825 2.74 ;
      RECT 0.605 2.06 1.825 2.265 ;
      RECT 0.605 0.33 0.775 2.265 ;
      RECT 2.565 0.82 2.815 1.49 ;
      RECT 0.605 0.82 2.815 0.99 ;
      RECT 0.605 0.33 0.785 0.99 ;
      RECT 0.38 0.33 0.785 0.66 ;
  END
END scs130lp_and4_0

MACRO scs130lp_and4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.495 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 0.805 1.345 1.475 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 0.805 1.825 1.475 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 1.345 2.355 1.76 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 0.255 3.275 3.075 ;
        RECT 2.69 0.255 3.275 1.015 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.25 -0.085 2.52 1.02 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.505 2.31 2.835 3.415 ;
        RECT 1.13 1.995 1.46 3.415 ;
        RECT 0.16 1.92 0.49 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.665 1.655 0.96 2.21 ;
      RECT 1.63 1.93 2.835 2.14 ;
      RECT 2.565 1.185 2.835 2.14 ;
      RECT 1.63 1.655 1.855 2.14 ;
      RECT 0.665 1.655 1.855 1.825 ;
      RECT 0.665 0.28 0.835 2.21 ;
      RECT 0.16 0.28 0.835 0.61 ;
  END
END scs130lp_and4_1

MACRO scs130lp_and4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.005 0.67 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.005 1.355 1.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.005 1.855 1.515 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 1.005 2.395 1.515 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 0.255 3.255 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.425 -0.085 3.715 1.105 ;
        RECT 2.36 -0.085 2.69 0.495 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.425 1.815 3.715 3.415 ;
        RECT 2.26 2.025 2.855 3.415 ;
        RECT 1.28 2.025 1.61 3.415 ;
        RECT 0.32 1.92 0.65 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.82 1.92 1.08 2.26 ;
      RECT 0.84 1.685 1.08 2.26 ;
      RECT 1.83 1.685 2.09 2.21 ;
      RECT 0.84 1.685 2.855 1.855 ;
      RECT 2.605 0.665 2.855 1.855 ;
      RECT 0.32 0.665 2.855 0.835 ;
      RECT 0.32 0.29 0.65 0.835 ;
  END
END scs130lp_and4_2

MACRO scs130lp_and4_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4_4 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.2 0.455 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.2 1.335 1.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.505 1.2 1.83 1.54 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 1.2 2.255 1.54 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.765 1.775 4.7 1.945 ;
        RECT 4.435 0.39 4.7 1.945 ;
        RECT 4.43 1.065 4.7 1.945 ;
        RECT 2.775 1.065 4.7 1.235 ;
        RECT 3.625 0.255 3.865 1.235 ;
        RECT 3.625 1.775 3.815 3.075 ;
        RECT 2.765 1.775 2.955 3.075 ;
        RECT 2.775 0.255 2.955 1.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.035 -0.085 4.265 0.895 ;
        RECT 3.125 -0.085 3.455 0.895 ;
        RECT 2.18 -0.085 2.51 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.985 2.115 4.315 3.415 ;
        RECT 3.125 2.115 3.455 3.415 ;
        RECT 2.18 2.105 2.51 3.415 ;
        RECT 1.185 2.105 1.515 3.415 ;
        RECT 0.25 1.92 0.58 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.685 1.755 2.01 3.075 ;
      RECT 0.75 1.755 1.015 3.075 ;
      RECT 0.75 1.755 2.595 1.925 ;
      RECT 2.425 0.86 2.595 1.925 ;
      RECT 2.425 1.415 4.26 1.585 ;
      RECT 0.31 0.86 2.595 1.03 ;
      RECT 0.31 0.36 0.5 1.03 ;
  END
END scs130lp_and4_4

MACRO scs130lp_and4_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4_lp 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.225 3.235 1.895 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.965 0.44 2.295 1.865 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 0.44 1.795 1.78 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 2.15 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 0.44 4.675 2.89 ;
        RECT 3.965 0.255 4.295 2.89 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.145 -0.085 3.475 0.715 ;
        RECT 0.585 -0.085 0.915 0.715 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.275 2.405 3.605 3.415 ;
        RECT 1.695 2.405 2.025 3.415 ;
        RECT 0.115 2.405 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.485 2.065 2.815 2.865 ;
      RECT 0.905 2.405 1.235 2.865 ;
      RECT 1.065 2.065 1.235 2.865 ;
      RECT 1.065 2.065 3.575 2.235 ;
      RECT 3.405 0.885 3.575 2.235 ;
      RECT 3.405 0.885 3.78 1.555 ;
      RECT 2.475 0.885 3.78 1.055 ;
      RECT 2.475 0.255 2.805 1.055 ;
  END
END scs130lp_and4_lp

MACRO scs130lp_and4_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4_lp2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.67 1.12 3.235 1.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.12 2.43 1.79 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.12 1.86 1.79 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.99 1.12 1.32 1.79 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.92 0.46 3.065 ;
        RECT 0.1 0.265 0.445 0.675 ;
        RECT 0.1 0.265 0.27 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 0.905 -0.085 1.235 0.59 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.895 2.025 3.225 3.415 ;
        RECT 1.755 2.32 2.085 3.415 ;
        RECT 0.66 2.32 0.99 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.365 1.97 2.695 3.065 ;
      RECT 1.225 1.97 1.555 3.065 ;
      RECT 0.64 1.97 2.695 2.14 ;
      RECT 0.64 0.77 0.81 2.14 ;
      RECT 0.45 0.94 0.81 1.61 ;
      RECT 2.615 0.265 2.945 0.94 ;
      RECT 0.64 0.77 2.945 0.94 ;
  END
END scs130lp_and4_lp2

MACRO scs130lp_and4_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.97 0.47 1.285 1.435 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.51 0.47 1.765 1.485 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.05 0.84 2.245 1.75 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 0.345 2.725 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.945 -0.085 2.275 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.085 2.065 2.295 3.415 ;
        RECT 1.225 2.065 1.435 3.415 ;
        RECT 0.365 2.065 0.575 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.655 1.715 1.865 3.045 ;
      RECT 0.79 1.715 1.005 2.265 ;
      RECT 0.62 1.715 1.865 1.885 ;
      RECT 0.62 0.33 0.79 1.885 ;
      RECT 0.285 0.33 0.79 0.66 ;
  END
END scs130lp_and4_m

MACRO scs130lp_and4b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4b_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.005 0.55 1.515 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.575 1.21 1.86 1.765 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 1.2 2.32 1.765 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.49 2.295 2.775 2.955 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 1.815 3.755 3.075 ;
        RECT 3.505 0.255 3.755 3.075 ;
        RECT 3.36 0.255 3.755 1.015 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.93 -0.085 3.19 1.015 ;
        RECT 2.555 -0.085 3.19 0.61 ;
        RECT 0.525 -0.085 0.855 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.945 1.815 3.265 3.415 ;
        RECT 2.9 1.815 3.265 2.125 ;
        RECT 1.585 1.935 2.32 3.415 ;
        RECT 0.6 2.035 0.93 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.49 1.185 2.73 2.125 ;
      RECT 1.11 1.795 1.405 2.125 ;
      RECT 1.235 0.255 1.405 2.125 ;
      RECT 2.49 1.185 3.335 1.515 ;
      RECT 2.49 0.86 2.67 2.125 ;
      RECT 1.235 0.86 2.67 1.03 ;
      RECT 1.235 0.255 1.515 1.03 ;
      RECT 1.045 0.255 1.515 0.485 ;
      RECT 0.15 1.695 0.43 2.21 ;
      RECT 0.15 1.695 0.93 1.865 ;
      RECT 0.76 0.655 0.93 1.865 ;
      RECT 0.76 0.655 1.065 1.445 ;
      RECT 0.095 0.655 1.065 0.825 ;
      RECT 0.095 0.29 0.355 0.825 ;
  END
END scs130lp_and4b_1

MACRO scs130lp_and4b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4b_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.815 0.425 1.485 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.575 1.21 1.835 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.175 2.35 1.75 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.52 1.175 2.89 1.54 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.6 0.86 3.78 1.88 ;
        RECT 3.475 1.71 3.7 3.075 ;
        RECT 3.41 0.255 3.66 1.04 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.95 -0.085 4.2 1.095 ;
        RECT 3.83 -0.085 4.2 0.69 ;
        RECT 2.91 -0.085 3.24 0.625 ;
        RECT 0.095 -0.085 0.425 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.885 2.05 4.2 3.415 ;
        RECT 3.95 1.815 4.2 3.415 ;
        RECT 2.88 2.05 3.305 3.415 ;
        RECT 1.575 1.92 2.305 3.415 ;
        RECT 0.655 2.035 0.985 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.52 1.71 2.71 2.25 ;
      RECT 1.155 0.795 1.405 2.25 ;
      RECT 2.52 1.71 3.24 1.88 ;
      RECT 3.07 0.795 3.24 1.88 ;
      RECT 3.07 1.21 3.43 1.54 ;
      RECT 1.075 0.795 3.24 1.005 ;
      RECT 0.225 1.695 0.475 2.25 ;
      RECT 0.225 1.695 0.795 1.865 ;
      RECT 0.595 0.255 0.795 1.865 ;
      RECT 0.595 0.255 1.255 0.595 ;
  END
END scs130lp_and4b_2

MACRO scs130lp_and4b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4b_4 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.38 0.815 2.19 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.94 1.335 4.645 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 1.345 3.77 1.75 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.965 1.345 3.265 1.75 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.855 2.455 2.26 ;
        RECT 0.985 1.075 2.455 1.245 ;
        RECT 2.265 0.255 2.455 1.245 ;
        RECT 1.365 0.255 1.595 1.245 ;
        RECT 0.985 1.075 1.165 2.26 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 2.7 -0.085 3.03 0.825 ;
        RECT 1.765 -0.085 2.095 0.905 ;
        RECT 0.985 -0.085 1.195 0.895 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.64 2.78 4.97 3.415 ;
        RECT 3.56 2.78 3.89 3.415 ;
        RECT 2.625 2.78 2.955 3.415 ;
        RECT 1.765 2.78 2.095 3.415 ;
        RECT 0.905 2.78 1.235 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.205 2.43 5.155 2.61 ;
      RECT 4.825 1.335 5.155 2.61 ;
      RECT 0.205 0.695 0.455 2.61 ;
      RECT 2.625 1.93 4.48 2.26 ;
      RECT 2.625 0.995 2.795 2.26 ;
      RECT 1.335 1.415 2.795 1.675 ;
      RECT 2.625 0.995 4.97 1.165 ;
      RECT 3.295 0.255 4.97 1.165 ;
  END
END scs130lp_and4b_4

MACRO scs130lp_and4b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4b_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 0.855 3.85 1.185 ;
        RECT 3.005 0.81 3.235 1.185 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.04 0.44 2.345 1.79 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 0.44 1.83 1.79 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.96 1.12 1.315 1.79 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 2.32 0.495 3.065 ;
        RECT 0.09 0.265 0.445 0.675 ;
        RECT 0.09 0.265 0.26 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.085 -0.085 3.415 0.63 ;
        RECT 0.905 -0.085 1.235 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.875 2.025 3.205 3.415 ;
        RECT 1.755 2.32 2.085 3.415 ;
        RECT 0.695 2.32 1.025 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.645 1.365 3.975 3.065 ;
      RECT 2.875 1.365 3.975 1.695 ;
      RECT 2.875 1.365 4.205 1.535 ;
      RECT 4.035 0.265 4.205 1.535 ;
      RECT 3.875 0.265 4.205 0.675 ;
      RECT 2.305 1.97 2.695 3.065 ;
      RECT 2.525 0.265 2.695 3.065 ;
      RECT 1.225 1.97 1.555 3.065 ;
      RECT 0.44 1.97 2.695 2.14 ;
      RECT 0.44 1.165 0.75 2.14 ;
      RECT 2.525 0.265 2.855 0.63 ;
  END
END scs130lp_and4b_lp

MACRO scs130lp_and4b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4b_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.055 0.55 1.565 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.47 1.895 1.485 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.47 2.435 1.565 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.805 0.84 3.205 1.565 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.45 0.47 3.685 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.85 -0.085 3.18 0.615 ;
        RECT 0.525 -0.085 0.855 0.525 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.99 2.095 3.2 3.415 ;
        RECT 1.96 2.155 2.29 3.415 ;
        RECT 1.11 2.095 1.32 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.48 2.855 2.81 3.025 ;
      RECT 2.48 1.745 2.69 3.025 ;
      RECT 1.57 1.745 1.78 2.295 ;
      RECT 1.22 1.745 2.69 1.915 ;
      RECT 1.22 0.475 1.41 1.915 ;
      RECT 0.68 1.745 0.89 2.295 ;
      RECT 0.84 0.705 1.01 1.915 ;
      RECT 0.155 0.705 1.01 0.875 ;
      RECT 0.155 0.385 0.345 0.875 ;
  END
END scs130lp_and4b_m

MACRO scs130lp_and4bb_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4bb_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.785 0.88 2.53 ;
        RECT 0.44 1.67 0.69 2.53 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.56 0.785 1.08 1.115 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.75 3.265 1.515 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.985 2.625 3.345 3.075 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.925 2.035 4.235 3.075 ;
        RECT 4.025 0.255 4.235 3.075 ;
        RECT 3.925 0.255 4.235 1.095 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.435 -0.085 3.755 1.095 ;
        RECT 0.56 -0.085 0.82 0.615 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.515 2.045 3.755 3.415 ;
        RECT 3.41 2.045 3.755 2.375 ;
        RECT 2.485 2.045 2.815 3.415 ;
        RECT 1.61 2.125 1.94 3.415 ;
        RECT 0.625 2.7 0.955 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.985 1.705 3.24 2.34 ;
      RECT 2.11 1.705 2.315 2.34 ;
      RECT 2.11 1.705 3.855 1.875 ;
      RECT 3.605 1.345 3.855 1.875 ;
      RECT 2.11 0.675 2.31 2.34 ;
      RECT 1.68 0.675 2.31 0.915 ;
      RECT 1.125 1.785 1.385 3.03 ;
      RECT 1.125 1.785 1.94 1.955 ;
      RECT 1.77 1.085 1.94 1.955 ;
      RECT 1.33 1.085 1.94 1.255 ;
      RECT 1.33 0.255 1.5 1.255 ;
      RECT 0.99 0.255 1.5 0.615 ;
      RECT 0.99 0.255 2.675 0.505 ;
      RECT 0.09 2.7 0.455 3.03 ;
      RECT 0.09 0.285 0.26 3.03 ;
      RECT 0.925 1.425 1.59 1.615 ;
      RECT 0.09 1.33 1.095 1.5 ;
      RECT 0.09 0.285 0.39 1.5 ;
  END
END scs130lp_and4bb_1

MACRO scs130lp_and4bb_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4bb_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.425 0.55 1.75 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.945 0.255 4.645 0.65 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.335 2.69 3.735 3.02 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.41 1.18 4.185 1.415 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.08 1.935 1.445 2.215 ;
        RECT 1.08 0.255 1.31 2.215 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.435 0.82 4.145 1.01 ;
        RECT 3.435 -0.085 3.775 1.01 ;
        RECT 1.48 -0.085 1.81 0.825 ;
        RECT 0.525 -0.085 0.91 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.905 2.12 4.185 3.415 ;
        RECT 2.985 2.275 3.315 2.52 ;
        RECT 2.985 2.275 3.155 3.415 ;
        RECT 1.545 2.725 2.22 3.415 ;
        RECT 1.955 2.135 2.22 3.415 ;
        RECT 0.685 2.725 1.015 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.355 0.82 4.685 2.45 ;
      RECT 2.79 1.585 4.685 1.765 ;
      RECT 2.79 1.245 3.12 1.765 ;
      RECT 3.485 1.935 3.735 2.45 ;
      RECT 2.39 1.935 2.815 2.45 ;
      RECT 2.39 1.935 3.735 2.105 ;
      RECT 2.39 0.67 2.56 2.45 ;
      RECT 1.48 0.995 1.75 1.615 ;
      RECT 1.48 0.995 2.56 1.175 ;
      RECT 2.125 0.67 2.56 1.175 ;
      RECT 0.73 2.385 1.785 2.555 ;
      RECT 1.615 1.795 1.785 2.555 ;
      RECT 0.16 1.92 0.9 2.385 ;
      RECT 1.615 1.795 2.22 1.965 ;
      RECT 1.96 1.345 2.22 1.965 ;
      RECT 0.73 1.075 0.9 2.555 ;
      RECT 0.095 1.075 0.9 1.245 ;
      RECT 0.095 0.71 0.355 1.245 ;
  END
END scs130lp_and4bb_2

MACRO scs130lp_and4bb_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4bb_4 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.69 1.425 6.14 1.76 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.47 0.855 2.12 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.48 1.21 3.9 1.79 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 1.21 3.31 1.795 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.075 2.515 1.245 ;
        RECT 2.325 0.255 2.515 1.245 ;
        RECT 1.115 1.815 2.505 2.145 ;
        RECT 1.425 0.255 1.655 1.245 ;
        RECT 1.115 1.075 1.295 2.145 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.385 -0.085 5.715 0.905 ;
        RECT 2.79 -0.085 3.12 0.7 ;
        RECT 1.825 -0.085 2.155 0.905 ;
        RECT 1.025 -0.085 1.255 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 4.77 2.815 5.1 3.415 ;
        RECT 3.75 2.815 4.08 3.415 ;
        RECT 2.765 2.815 3.095 3.415 ;
        RECT 1.825 2.815 2.155 3.415 ;
        RECT 0.965 2.815 1.295 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.34 1.93 5.64 2.26 ;
      RECT 5.34 1.075 5.51 2.26 ;
      RECT 4.645 1.075 4.975 1.445 ;
      RECT 4.645 1.075 6.145 1.245 ;
      RECT 5.885 0.695 6.145 1.245 ;
      RECT 2.685 1.965 4.61 2.295 ;
      RECT 2.685 0.87 2.855 2.295 ;
      RECT 1.465 1.415 2.855 1.645 ;
      RECT 2.685 0.87 4.405 1.04 ;
      RECT 3.46 0.255 5.1 0.905 ;
      RECT 0.205 2.465 4.96 2.645 ;
      RECT 4.79 1.615 4.96 2.645 ;
      RECT 0.205 0.7 0.455 2.645 ;
      RECT 4.105 1.615 4.96 1.785 ;
      RECT 4.105 1.345 4.445 1.785 ;
  END
END scs130lp_and4bb_4

MACRO scs130lp_and4bb_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4bb_lp 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.785 1.315 1.455 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.125 1.89 1.455 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.37 1.12 3.715 1.79 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.94 1.12 4.27 1.79 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.8 1.92 5.19 3.065 ;
        RECT 5.02 0.265 5.19 3.065 ;
        RECT 4.815 0.265 5.19 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 3.885 -0.085 4.215 0.59 ;
        RECT 0.905 -0.085 1.235 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.165 2.32 4.495 3.415 ;
        RECT 3.025 2.685 3.355 3.415 ;
        RECT 1.965 2.335 2.295 3.415 ;
        RECT 0.645 1.985 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.635 1.97 3.965 3.065 ;
      RECT 2.495 2.335 2.825 3.065 ;
      RECT 2.495 2.335 3.965 2.505 ;
      RECT 3.635 1.97 4.62 2.14 ;
      RECT 4.45 0.77 4.62 2.14 ;
      RECT 4.45 0.94 4.84 1.61 ;
      RECT 3.31 0.77 4.62 0.94 ;
      RECT 3.31 0.265 3.48 0.94 ;
      RECT 2.285 0.265 3.48 0.595 ;
      RECT 1.435 1.985 1.765 3.065 ;
      RECT 1.435 1.985 2.97 2.155 ;
      RECT 2.8 0.775 2.97 2.155 ;
      RECT 2.8 1.215 3.13 1.885 ;
      RECT 1.725 0.775 2.97 0.945 ;
      RECT 1.725 0.265 2.055 0.945 ;
      RECT 0.115 0.265 0.445 3.025 ;
      RECT 0.115 1.635 2.56 1.805 ;
      RECT 2.23 1.135 2.56 1.805 ;
  END
END scs130lp_and4bb_lp

MACRO scs130lp_and4bb_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_and4bb_m 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.475 0.805 0.805 1.475 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 0.805 1.285 1.475 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.975 1.405 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.95 3.335 2.12 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.73 2.655 4.165 2.985 ;
        RECT 3.975 0.47 4.165 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.505 -0.085 3.715 0.935 ;
        RECT 0.72 -0.085 0.93 0.585 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.22 2.845 3.55 3.415 ;
        RECT 2.4 2.785 2.61 3.415 ;
        RECT 1.54 2.785 1.75 3.415 ;
        RECT 0.72 2.095 0.93 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.83 2.435 3.04 2.985 ;
      RECT 1.97 2.435 2.18 2.985 ;
      RECT 1.97 2.435 3.04 2.605 ;
      RECT 2.655 1.585 2.825 2.605 ;
      RECT 3.625 1.585 3.795 2.255 ;
      RECT 2.655 1.585 3.795 1.755 ;
      RECT 3.155 0.645 3.325 1.755 ;
      RECT 1.68 0.645 3.325 0.975 ;
      RECT 1.15 0.265 1.36 0.595 ;
      RECT 1.15 0.265 2.615 0.435 ;
      RECT 1.15 2.005 1.36 2.335 ;
      RECT 1.15 2.005 2.435 2.175 ;
      RECT 2.105 1.615 2.435 2.175 ;
      RECT 0.125 1.655 0.5 2.295 ;
      RECT 0.125 1.655 1.785 1.825 ;
      RECT 1.615 1.155 1.785 1.825 ;
      RECT 0.125 0.295 0.295 2.295 ;
      RECT 0.125 0.295 0.5 0.625 ;
  END
END scs130lp_and4bb_m

MACRO scs130lp_buf_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_0 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.89 1.15 1.345 1.885 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 2.395 0.4 3.075 ;
        RECT 0.09 0.285 0.39 0.615 ;
        RECT 0.09 1.605 0.34 3.075 ;
        RECT 0.09 0.285 0.26 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.56 -0.085 0.89 0.615 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.57 2.395 0.825 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.995 2.055 1.345 3.075 ;
      RECT 0.51 2.055 1.345 2.225 ;
      RECT 0.51 0.785 0.68 2.225 ;
      RECT 0.43 0.785 0.68 1.455 ;
      RECT 0.43 0.785 1.345 0.97 ;
      RECT 1.06 0.3 1.345 0.97 ;
  END
END scs130lp_buf_0

MACRO scs130lp_buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 1.19 1.355 1.435 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.865 0.355 3.075 ;
        RECT 0.085 0.255 0.355 1.03 ;
        RECT 0.085 0.255 0.26 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.525 -0.085 0.855 0.68 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.525 1.945 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.025 1.605 1.345 2.485 ;
      RECT 0.505 1.605 1.345 1.775 ;
      RECT 0.43 1.185 0.695 1.705 ;
      RECT 0.525 0.85 0.695 1.775 ;
      RECT 0.525 0.85 1.345 1.02 ;
      RECT 1.025 0.69 1.345 1.02 ;
  END
END scs130lp_buf_1

MACRO scs130lp_buf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_16 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.89 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.365 1.385 2.735 1.585 ;
        RECT 1.905 1.205 2.255 1.585 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    ANTENNADIFFAREA 4.704 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 3.225 1.92 9.535 2.15 ;
      LAYER li ;
        RECT 9.26 0.255 9.52 3.075 ;
        RECT 8.4 0.255 8.66 3.075 ;
        RECT 7.54 0.255 7.8 3.075 ;
        RECT 6.68 0.255 6.94 3.075 ;
        RECT 5.82 0.255 6.08 3.075 ;
        RECT 4.96 0.255 5.22 3.075 ;
        RECT 4.1 0.255 4.36 3.075 ;
        RECT 3.265 0.255 3.5 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.69 -0.085 9.985 1.075 ;
        RECT 8.83 -0.085 9.09 1.075 ;
        RECT 7.97 -0.085 8.23 1.075 ;
        RECT 7.11 -0.085 7.37 1.075 ;
        RECT 6.25 -0.085 6.51 1.075 ;
        RECT 5.39 -0.085 5.65 1.075 ;
        RECT 4.53 -0.085 4.79 1.075 ;
        RECT 3.67 -0.085 3.93 1.075 ;
        RECT 2.81 -0.085 3.095 0.875 ;
        RECT 1.915 -0.085 2.245 0.695 ;
        RECT 1.09 -0.085 1.36 0.875 ;
        RECT 0.195 -0.085 0.49 1.075 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.69 1.92 9.985 3.415 ;
        RECT 8.83 1.92 9.09 3.415 ;
        RECT 7.97 1.92 8.23 3.415 ;
        RECT 7.11 1.92 7.37 3.415 ;
        RECT 6.25 1.92 6.51 3.415 ;
        RECT 5.39 1.92 5.65 3.415 ;
        RECT 4.53 1.92 4.79 3.415 ;
        RECT 3.67 1.92 3.93 3.415 ;
        RECT 2.81 2.095 3.095 3.415 ;
        RECT 1.95 2.095 2.21 3.415 ;
        RECT 1.09 2.095 1.35 3.415 ;
        RECT 0.195 1.815 0.49 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 2.855 1.55 9.105 1.78 ;
    LAYER li ;
      RECT 2.38 1.755 2.64 3.075 ;
      RECT 1.52 1.755 1.78 3.075 ;
      RECT 0.66 1.755 0.92 3.075 ;
      RECT 0.66 1.755 3.095 1.925 ;
      RECT 2.905 1.045 3.095 1.925 ;
      RECT 2.425 1.045 3.095 1.215 ;
      RECT 0.66 1.045 1.735 1.215 ;
      RECT 1.53 0.425 1.735 1.215 ;
      RECT 2.425 0.425 2.64 1.215 ;
      RECT 0.66 0.425 0.92 1.215 ;
      RECT 1.53 0.865 2.64 1.035 ;
      RECT 2.415 0.425 2.64 1.035 ;
      RECT 1.53 0.425 1.745 1.035 ;
      RECT 8.83 1.325 9.09 1.75 ;
      RECT 7.97 1.325 8.23 1.75 ;
      RECT 7.11 1.325 7.37 1.75 ;
      RECT 6.25 1.325 6.51 1.75 ;
      RECT 5.39 1.325 5.65 1.75 ;
      RECT 4.53 1.325 4.79 1.75 ;
      RECT 3.67 1.325 3.93 1.75 ;
  END
END scs130lp_buf_16

MACRO scs130lp_buf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 1.185 1.785 1.515 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.61 2.045 0.875 3.055 ;
        RECT 0.61 0.255 0.835 3.055 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.005 -0.085 1.785 1.015 ;
        RECT 0.145 -0.085 0.44 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.045 2.025 1.785 3.415 ;
        RECT 0.245 2.105 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.955 0.7 2.215 2.485 ;
      RECT 1.005 1.685 2.215 1.855 ;
      RECT 1.005 1.345 1.275 1.855 ;
  END
END scs130lp_buf_2

MACRO scs130lp_buf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_4 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.39 1.2 2.785 1.54 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.665 1.775 1.855 3.075 ;
        RECT 0.095 1.075 1.855 1.245 ;
        RECT 1.665 0.255 1.855 1.245 ;
        RECT 0.095 1.775 1.855 1.945 ;
        RECT 0.805 1.775 0.995 3.075 ;
        RECT 0.805 0.255 0.995 1.245 ;
        RECT 0.095 1.075 0.51 1.945 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.025 -0.085 2.355 0.69 ;
        RECT 1.165 -0.085 1.495 0.905 ;
        RECT 0.305 -0.085 0.635 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.025 2.095 2.355 3.415 ;
        RECT 1.165 2.115 1.495 3.415 ;
        RECT 0.305 2.115 0.635 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.525 1.755 2.785 3.075 ;
      RECT 2.025 1.755 2.785 1.925 ;
      RECT 2.025 0.86 2.22 1.925 ;
      RECT 0.7 1.415 2.22 1.605 ;
      RECT 2.025 0.86 2.785 1.03 ;
      RECT 2.525 0.255 2.785 1.03 ;
  END
END scs130lp_buf_4

MACRO scs130lp_buf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_8 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.945 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.385 1.345 1.575 ;
        RECT 0.095 1.18 0.88 1.575 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.865 1.745 5.19 1.925 ;
        RECT 4.91 1.045 5.19 1.925 ;
        RECT 1.865 1.045 5.19 1.225 ;
        RECT 4.43 1.745 4.69 2.98 ;
        RECT 4.43 0.305 4.685 1.225 ;
        RECT 3.57 1.745 3.83 2.98 ;
        RECT 3.57 0.305 3.83 1.225 ;
        RECT 2.705 1.745 2.975 2.98 ;
        RECT 2.71 0.305 2.965 1.225 ;
        RECT 1.865 0.305 2.11 1.225 ;
        RECT 1.865 1.745 2.105 2.98 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.855 -0.085 5.155 0.875 ;
        RECT 4 -0.085 4.26 0.875 ;
        RECT 3.135 -0.085 3.4 0.875 ;
        RECT 2.28 -0.085 2.54 0.875 ;
        RECT 1.42 -0.085 1.695 0.875 ;
        RECT 0.56 -0.085 0.82 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.86 2.095 5.095 3.415 ;
        RECT 4 2.095 4.26 3.415 ;
        RECT 3.145 2.095 3.4 3.415 ;
        RECT 2.275 2.095 2.535 3.415 ;
        RECT 1.42 2.095 1.695 3.415 ;
        RECT 0.56 2.095 0.82 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.99 1.745 1.25 2.98 ;
      RECT 0.095 1.745 0.39 2.98 ;
      RECT 0.095 1.745 1.695 1.925 ;
      RECT 1.525 1.045 1.695 1.925 ;
      RECT 1.525 1.395 4.74 1.575 ;
      RECT 1.05 1.045 1.695 1.215 ;
      RECT 1.05 0.305 1.25 1.215 ;
      RECT 0.095 0.84 1.25 1.01 ;
      RECT 0.99 0.305 1.25 1.01 ;
      RECT 0.095 0.305 0.39 1.01 ;
  END
END scs130lp_buf_8

MACRO scs130lp_buf_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 0.44 1.795 1.485 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.23 1.835 0.56 3.055 ;
        RECT 0.125 0.265 0.495 2.89 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.955 -0.085 1.285 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.76 2.015 1.09 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.535 1.665 1.865 3.055 ;
      RECT 0.74 1.665 2.225 1.835 ;
      RECT 1.975 0.265 2.225 1.835 ;
      RECT 0.74 1.165 1.07 1.835 ;
  END
END scs130lp_buf_lp

MACRO scs130lp_buf_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buf_m 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 0.875 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.46 0.365 2.96 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.585 -0.085 0.795 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.585 2.76 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.015 1.93 1.225 2.96 ;
      RECT 1.055 0.33 1.225 2.96 ;
      RECT 0.545 1.93 1.225 2.1 ;
      RECT 1.015 0.33 1.225 0.66 ;
  END
END scs130lp_buf_m

MACRO scs130lp_bufbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufbuf_16 0 0 ;
  SIZE 12.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.355 0.485 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    ANTENNADIFFAREA 4.704 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 5.625 1.92 11.935 2.15 ;
      LAYER li ;
        RECT 11.66 0.255 11.92 3.075 ;
        RECT 10.8 0.255 11.06 3.075 ;
        RECT 9.94 0.255 10.2 3.075 ;
        RECT 9.08 0.255 9.34 3.075 ;
        RECT 8.22 0.255 8.48 3.075 ;
        RECT 7.36 0.255 7.62 3.075 ;
        RECT 6.5 0.255 6.76 3.075 ;
        RECT 5.665 0.255 5.9 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.48 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.48 0.085 ;
        RECT 12.09 -0.085 12.385 1.075 ;
        RECT 11.23 -0.085 11.49 1.075 ;
        RECT 10.37 -0.085 10.63 1.075 ;
        RECT 9.51 -0.085 9.77 1.075 ;
        RECT 8.65 -0.085 8.91 1.075 ;
        RECT 7.79 -0.085 8.05 1.075 ;
        RECT 6.93 -0.085 7.19 1.075 ;
        RECT 6.07 -0.085 6.33 1.075 ;
        RECT 5.21 -0.085 5.47 0.875 ;
        RECT 4.35 -0.085 4.61 0.875 ;
        RECT 3.455 -0.085 3.75 0.875 ;
        RECT 2.595 -0.085 2.885 0.895 ;
        RECT 1.385 -0.085 1.715 0.895 ;
        RECT 0.525 -0.085 0.855 0.845 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.48 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.48 3.415 ;
        RECT 12.09 1.925 12.385 3.415 ;
        RECT 11.23 1.925 11.49 3.415 ;
        RECT 10.37 1.925 10.63 3.415 ;
        RECT 9.51 1.925 9.77 3.415 ;
        RECT 8.65 1.925 8.91 3.415 ;
        RECT 7.79 1.925 8.05 3.415 ;
        RECT 6.93 1.925 7.19 3.415 ;
        RECT 6.07 1.925 6.33 3.415 ;
        RECT 5.21 2.095 5.47 3.415 ;
        RECT 4.35 2.095 4.61 3.415 ;
        RECT 3.49 2.095 3.75 3.415 ;
        RECT 2.595 2.1 2.925 3.415 ;
        RECT 1.385 2.115 1.715 3.415 ;
        RECT 0.56 2.26 0.82 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 5.255 1.55 11.505 1.78 ;
    LAYER li ;
      RECT 4.78 1.745 5.04 3.075 ;
      RECT 3.92 1.745 4.18 3.075 ;
      RECT 3.095 1.745 3.32 3.075 ;
      RECT 3.095 1.745 5.495 1.925 ;
      RECT 5.305 1.045 5.495 1.925 ;
      RECT 3.055 1.045 5.495 1.215 ;
      RECT 4.78 0.255 5.04 1.215 ;
      RECT 3.92 0.255 4.18 1.215 ;
      RECT 3.055 0.255 3.285 1.215 ;
      RECT 1.885 1.76 2.145 3.075 ;
      RECT 1.005 1.76 1.215 3.075 ;
      RECT 1.005 1.76 2.145 1.945 ;
      RECT 1.005 1.76 2.52 1.93 ;
      RECT 2.35 1.065 2.52 1.93 ;
      RECT 2.35 1.385 5.135 1.575 ;
      RECT 2.35 1.065 2.855 1.575 ;
      RECT 1.025 1.065 2.855 1.235 ;
      RECT 1.885 0.255 2.145 1.235 ;
      RECT 1.025 0.255 1.215 1.235 ;
      RECT 0.095 1.92 0.39 3.075 ;
      RECT 0.095 1.92 0.835 2.09 ;
      RECT 0.665 1.015 0.835 2.09 ;
      RECT 0.665 1.405 2.18 1.59 ;
      RECT 0.095 1.015 0.835 1.185 ;
      RECT 0.095 0.255 0.355 1.185 ;
      RECT 11.23 1.315 11.49 1.755 ;
      RECT 10.37 1.315 10.63 1.755 ;
      RECT 9.51 1.315 9.77 1.755 ;
      RECT 8.65 1.315 8.91 1.755 ;
      RECT 7.79 1.315 8.05 1.755 ;
      RECT 6.93 1.315 7.19 1.755 ;
      RECT 6.07 1.315 6.33 1.755 ;
  END
END scs130lp_bufbuf_16

MACRO scs130lp_bufbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufbuf_8 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.65 1.405 7.115 1.755 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.44 1.755 3.665 3.075 ;
        RECT 0.085 1.055 3.665 1.225 ;
        RECT 3.475 0.29 3.665 1.225 ;
        RECT 0.085 1.755 3.665 1.925 ;
        RECT 2.58 1.755 2.84 3.075 ;
        RECT 2.615 0.29 2.805 1.225 ;
        RECT 1.72 1.755 1.98 3.075 ;
        RECT 1.755 0.29 1.945 1.225 ;
        RECT 0.86 1.755 1.12 3.075 ;
        RECT 0.895 0.29 1.085 1.225 ;
        RECT 0.085 1.055 0.405 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 6.21 -0.085 6.54 0.895 ;
        RECT 4.74 -0.085 5.07 0.885 ;
        RECT 3.835 -0.085 4.19 0.885 ;
        RECT 2.975 -0.085 3.305 0.885 ;
        RECT 2.115 -0.085 2.445 0.885 ;
        RECT 1.255 -0.085 1.585 0.885 ;
        RECT 0.395 -0.085 0.725 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.25 2.37 6.58 3.415 ;
        RECT 4.78 2.095 5.04 3.415 ;
        RECT 3.835 2.095 4.165 3.415 ;
        RECT 3.01 2.105 3.27 3.415 ;
        RECT 2.15 2.105 2.41 3.415 ;
        RECT 1.29 2.105 1.55 3.415 ;
        RECT 0.395 2.105 0.69 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.24 1.925 7.105 2.2 ;
      RECT 6.24 1.065 6.44 2.2 ;
      RECT 6.19 1.065 6.44 1.525 ;
      RECT 6.19 1.065 7.105 1.235 ;
      RECT 6.775 0.665 7.105 1.235 ;
      RECT 5.84 1.815 6.07 2.825 ;
      RECT 5.84 0.435 6.02 2.825 ;
      RECT 4.185 1.395 6.02 1.585 ;
      RECT 5.76 0.435 6.02 1.585 ;
      RECT 5.21 1.755 5.5 3.075 ;
      RECT 4.335 1.755 4.61 3.075 ;
      RECT 3.835 1.755 5.5 1.925 ;
      RECT 3.835 1.055 4.005 1.925 ;
      RECT 0.585 1.395 4.005 1.585 ;
      RECT 3.835 1.055 5.5 1.225 ;
      RECT 5.24 0.29 5.5 1.225 ;
      RECT 4.36 0.29 4.57 1.225 ;
  END
END scs130lp_bufbuf_8

MACRO scs130lp_bufinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufinv_16 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.945 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.415 1.57 1.76 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    ANTENNADIFFAREA 4.704 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 4.64 1.92 10.95 2.15 ;
      LAYER li ;
        RECT 10.675 0.315 10.935 3.025 ;
        RECT 9.815 0.315 10.075 3.025 ;
        RECT 8.955 0.315 9.215 3.025 ;
        RECT 8.095 0.315 8.355 3.025 ;
        RECT 7.235 0.315 7.495 3.025 ;
        RECT 6.375 0.315 6.635 3.025 ;
        RECT 5.515 0.315 5.775 3.025 ;
        RECT 4.69 0.315 4.915 3.025 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.52 0.085 ;
        RECT 11.105 -0.085 11.4 1.08 ;
        RECT 10.245 -0.085 10.505 1.08 ;
        RECT 9.385 -0.085 9.645 1.08 ;
        RECT 8.525 -0.085 8.785 1.08 ;
        RECT 7.665 -0.085 7.925 1.08 ;
        RECT 6.805 -0.085 7.065 1.08 ;
        RECT 5.945 -0.085 6.205 1.08 ;
        RECT 5.085 -0.085 5.345 1.08 ;
        RECT 4.225 -0.085 4.485 0.885 ;
        RECT 3.365 -0.085 3.625 0.885 ;
        RECT 2.505 -0.085 2.765 0.885 ;
        RECT 1.6 -0.085 1.87 0.905 ;
        RECT 0.74 -0.085 1 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.52 3.415 ;
        RECT 11.105 1.955 11.4 3.415 ;
        RECT 10.245 1.955 10.505 3.415 ;
        RECT 9.385 1.955 9.645 3.415 ;
        RECT 8.525 1.955 8.785 3.415 ;
        RECT 7.665 1.955 7.925 3.415 ;
        RECT 6.805 1.955 7.065 3.415 ;
        RECT 5.945 1.955 6.205 3.415 ;
        RECT 5.085 1.955 5.345 3.415 ;
        RECT 4.225 2.105 4.485 3.415 ;
        RECT 3.365 2.105 3.625 3.415 ;
        RECT 2.505 2.105 2.765 3.415 ;
        RECT 1.6 2.27 1.905 3.415 ;
        RECT 0.74 2.27 1 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 4.29 1.55 10.52 1.78 ;
    LAYER li ;
      RECT 3.795 1.755 4.055 3.025 ;
      RECT 2.935 1.755 3.195 3.025 ;
      RECT 2.09 1.755 2.335 3.025 ;
      RECT 2.09 1.755 4.52 1.925 ;
      RECT 4.34 1.055 4.52 1.925 ;
      RECT 2.09 1.055 4.52 1.225 ;
      RECT 3.795 0.315 4.055 1.225 ;
      RECT 2.935 0.315 3.195 1.225 ;
      RECT 2.09 0.315 2.335 1.225 ;
      RECT 1.17 1.93 1.43 3.025 ;
      RECT 0.275 1.93 0.57 3.025 ;
      RECT 0.275 1.93 1.92 2.1 ;
      RECT 1.75 1.075 1.92 2.1 ;
      RECT 1.75 1.395 4.17 1.585 ;
      RECT 0.275 1.075 1.92 1.245 ;
      RECT 1.17 0.315 1.43 1.245 ;
      RECT 0.275 0.315 0.57 1.245 ;
      RECT 10.245 1.345 10.505 1.785 ;
      RECT 9.385 1.345 9.645 1.785 ;
      RECT 8.525 1.345 8.785 1.785 ;
      RECT 7.665 1.345 7.925 1.785 ;
      RECT 6.805 1.345 7.065 1.785 ;
      RECT 5.945 1.345 6.205 1.785 ;
      RECT 5.085 1.345 5.345 1.785 ;
  END
END scs130lp_bufinv_16

MACRO scs130lp_bufinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufinv_8 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.75 1.21 6.155 1.8 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.15 1.755 3.41 3.055 ;
        RECT 3.15 0.255 3.41 1.225 ;
        RECT 0.095 1.755 3.41 1.925 ;
        RECT 0.57 1.055 3.41 1.225 ;
        RECT 2.29 1.755 2.55 3.055 ;
        RECT 2.29 0.255 2.55 1.225 ;
        RECT 1.43 1.755 1.69 3.055 ;
        RECT 1.43 0.255 1.69 1.225 ;
        RECT 0.57 1.755 0.83 3.055 ;
        RECT 0.57 0.255 0.83 1.225 ;
        RECT 0.095 1.16 0.815 1.925 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.365 -0.085 5.695 0.7 ;
        RECT 4.505 -0.085 4.835 0.885 ;
        RECT 3.58 -0.085 3.86 1.07 ;
        RECT 2.72 -0.085 2.98 0.885 ;
        RECT 1.86 -0.085 2.12 0.885 ;
        RECT 1 -0.085 1.26 0.885 ;
        RECT 0.105 -0.085 0.4 0.99 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.365 2.31 5.695 3.415 ;
        RECT 4.545 2.095 4.8 3.415 ;
        RECT 3.58 1.84 3.87 3.415 ;
        RECT 2.72 2.095 2.98 3.415 ;
        RECT 1.86 2.095 2.12 3.415 ;
        RECT 1 2.095 1.26 3.415 ;
        RECT 0.105 2.095 0.4 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.865 1.97 6.125 3.055 ;
      RECT 5.385 1.97 6.125 2.14 ;
      RECT 5.385 0.87 5.555 2.14 ;
      RECT 4.38 1.395 5.555 1.585 ;
      RECT 5.385 0.87 6.145 1.04 ;
      RECT 5.865 0.255 6.145 1.04 ;
      RECT 4.97 1.755 5.195 3.055 ;
      RECT 4.04 1.755 4.375 3.055 ;
      RECT 4.04 1.755 5.195 1.925 ;
      RECT 4.04 0.255 4.21 3.055 ;
      RECT 0.985 1.395 4.21 1.585 ;
      RECT 4.03 0.255 4.21 1.585 ;
      RECT 4.03 1.055 5.195 1.225 ;
      RECT 5.005 0.255 5.195 1.225 ;
      RECT 4.03 0.255 4.335 1.225 ;
  END
END scs130lp_bufinv_8

MACRO scs130lp_bufkapwr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufkapwr_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.345 1.015 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.3 0.43 0.635 ;
        RECT 0.085 1.525 0.395 3.075 ;
        RECT 0.085 0.3 0.255 3.075 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 1.37 2.945 ;
      LAYER li ;
        RECT 0.565 1.92 0.825 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.6 -0.085 0.875 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.995 1.92 1.355 3.075 ;
      RECT 1.185 0.3 1.355 3.075 ;
      RECT 0.425 0.805 1.355 1.135 ;
      RECT 1.045 0.3 1.355 1.135 ;
  END
END scs130lp_bufkapwr_1

MACRO scs130lp_bufkapwr_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufkapwr_2 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.425 0.775 0.875 1.105 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.725 1.815 1.895 ;
        RECT 1.385 0.78 1.815 1.895 ;
        RECT 1.045 0.78 1.815 1.105 ;
        RECT 1.045 1.725 1.305 3.045 ;
        RECT 1.045 0.265 1.305 1.105 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 1.85 2.945 ;
      LAYER li ;
        RECT 1.475 2.065 1.73 3.075 ;
        RECT 0.565 1.875 0.875 3.045 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.475 -0.085 1.73 0.61 ;
        RECT 0.555 -0.085 0.83 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.275 0.395 3.045 ;
      RECT 0.085 1.275 1.215 1.535 ;
      RECT 0.085 0.265 0.255 3.045 ;
      RECT 0.085 0.265 0.385 0.605 ;
  END
END scs130lp_bufkapwr_2

MACRO scs130lp_bufkapwr_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufkapwr_4 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.425 0.775 0.805 1.105 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9408 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.725 2.765 1.895 ;
        RECT 2.255 0.775 2.765 1.895 ;
        RECT 1.045 0.775 2.765 1.025 ;
        RECT 1.905 1.725 2.165 3.06 ;
        RECT 1.905 0.275 2.165 1.025 ;
        RECT 1.045 1.725 1.305 3.06 ;
        RECT 1.045 0.275 1.305 1.025 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 2.81 2.945 ;
      LAYER li ;
        RECT 2.335 2.065 2.62 3.075 ;
        RECT 1.475 2.065 1.73 3.075 ;
        RECT 0.565 1.875 0.875 3.06 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.335 -0.085 2.615 0.605 ;
        RECT 1.475 -0.085 1.73 0.605 ;
        RECT 0.555 -0.085 0.83 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.275 0.395 3.06 ;
      RECT 0.085 1.275 2.085 1.535 ;
      RECT 1.075 1.205 2.085 1.535 ;
      RECT 0.085 0.275 0.255 3.06 ;
      RECT 0.085 0.275 0.385 0.605 ;
  END
END scs130lp_bufkapwr_4

MACRO scs130lp_bufkapwr_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bufkapwr_8 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.4 1.57 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8816 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.42 1.655 4.73 1.895 ;
        RECT 3.76 0.735 4.73 1.895 ;
        RECT 4 0.28 4.26 3.075 ;
        RECT 1.42 0.735 4.73 0.975 ;
        RECT 3.14 1.655 3.4 3.075 ;
        RECT 3.14 0.28 3.4 0.975 ;
        RECT 2.28 1.655 2.54 3.075 ;
        RECT 2.28 0.28 2.54 0.975 ;
        RECT 1.42 1.655 1.68 3.075 ;
        RECT 1.42 0.28 1.68 0.975 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 5.21 2.945 ;
      LAYER li ;
        RECT 4.43 2.065 4.725 3.075 ;
        RECT 3.57 2.065 3.83 3.075 ;
        RECT 2.71 2.065 2.97 3.075 ;
        RECT 1.85 2.065 2.11 3.075 ;
        RECT 0.99 1.875 1.25 3.055 ;
        RECT 0.095 1.875 0.39 3.055 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.43 -0.085 4.73 0.565 ;
        RECT 3.57 -0.085 3.83 0.565 ;
        RECT 2.71 -0.085 2.97 0.565 ;
        RECT 1.85 -0.085 2.11 0.565 ;
        RECT 0.99 -0.085 1.25 0.61 ;
        RECT 0.145 -0.085 0.39 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.57 0.265 0.82 3.075 ;
      RECT 0.57 1.155 3.59 1.485 ;
  END
END scs130lp_bufkapwr_8

MACRO scs130lp_buflp_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buflp_0 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.55 0.935 2.89 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3021 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.8 0.44 2.275 2.89 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.98 -0.085 1.31 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.12 2.21 1.45 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.16 0.58 0.435 2.89 ;
      RECT 1.245 1.21 1.575 1.88 ;
      RECT 0.16 1.21 1.575 1.38 ;
      RECT 0.16 0.58 0.49 1.38 ;
  END
END scs130lp_buflp_0

MACRO scs130lp_buflp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buflp_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.445 1.185 1.795 2.89 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.255 0.455 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.945 -0.085 1.275 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.945 1.815 1.275 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.985 0.635 2.235 2.675 ;
      RECT 0.82 0.845 1.15 1.515 ;
      RECT 0.82 0.845 2.235 1.015 ;
      RECT 1.905 0.635 2.235 1.015 ;
  END
END scs130lp_buflp_1

MACRO scs130lp_buflp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buflp_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 1.055 2.805 2.89 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6468 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.595 1.445 1.095 ;
        RECT 1.045 1.55 1.375 2.735 ;
        RECT 1.115 0.595 1.375 2.735 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.115 -0.085 2.445 0.545 ;
        RECT 0.115 -0.085 0.445 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.975 1.815 2.305 3.415 ;
        RECT 0.115 1.815 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.99 0.255 3.245 2.545 ;
      RECT 1.825 1.265 2.285 1.595 ;
      RECT 2.115 0.715 2.285 1.595 ;
      RECT 2.115 0.715 3.245 0.885 ;
      RECT 2.915 0.255 3.245 0.885 ;
      RECT 1.615 0.255 1.945 1.095 ;
      RECT 0.615 0.255 0.945 1.095 ;
      RECT 0.615 0.255 1.945 0.425 ;
      RECT 0.615 2.905 1.805 3.075 ;
      RECT 1.555 1.815 1.805 3.075 ;
      RECT 0.615 1.815 0.865 3.075 ;
  END
END scs130lp_buflp_2

MACRO scs130lp_buflp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buflp_4 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 1.18 4.43 1.515 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3524 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.815 3.235 2.735 ;
        RECT 0.125 0.975 2.945 1.145 ;
        RECT 2.775 0.595 2.945 1.145 ;
        RECT 0.185 1.815 3.235 1.985 ;
        RECT 1.905 1.815 2.235 2.735 ;
        RECT 1.835 0.595 2.085 1.145 ;
        RECT 0.185 0.975 0.355 1.985 ;
        RECT 0.125 0.975 0.355 1.78 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 3.625 -0.085 3.955 0.67 ;
        RECT 0.975 -0.085 1.305 0.465 ;
        RECT 0.115 -0.085 0.365 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 3.905 1.815 4.235 3.415 ;
        RECT 1.055 2.495 1.225 3.415 ;
        RECT 0.115 2.155 0.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.795 0.255 5.125 3.075 ;
      RECT 0.745 1.315 3.795 1.645 ;
      RECT 3.625 0.84 3.795 1.645 ;
      RECT 3.625 0.84 5.125 1.01 ;
      RECT 1.405 2.905 3.735 3.075 ;
      RECT 3.405 1.815 3.735 3.075 ;
      RECT 0.545 2.155 0.875 3.075 ;
      RECT 2.405 2.155 2.735 3.075 ;
      RECT 1.405 2.155 1.735 3.075 ;
      RECT 0.545 2.155 1.735 2.325 ;
      RECT 3.125 0.255 3.455 1.095 ;
      RECT 2.265 0.255 2.595 0.805 ;
      RECT 0.545 0.635 1.655 0.805 ;
      RECT 1.485 0.255 1.655 0.805 ;
      RECT 0.545 0.255 0.795 0.805 ;
      RECT 1.485 0.255 3.455 0.425 ;
  END
END scs130lp_buflp_4

MACRO scs130lp_buflp_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buflp_8 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.89 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.535 1.185 2.565 1.515 ;
        RECT 0.535 1.18 2.255 1.515 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8224 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.235 1.765 10.435 1.935 ;
        RECT 9.995 0.925 10.435 1.935 ;
        RECT 6.405 0.925 10.435 1.095 ;
        RECT 9.235 1.765 9.565 2.735 ;
        RECT 9.185 0.595 9.515 1.095 ;
        RECT 8.235 1.765 8.565 2.735 ;
        RECT 8.185 0.595 8.515 1.095 ;
        RECT 7.235 1.765 7.565 2.735 ;
        RECT 7.265 0.595 7.515 1.095 ;
        RECT 6.405 0.595 6.575 1.095 ;
        RECT 6.235 1.765 6.565 2.735 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 10.115 -0.085 10.445 0.755 ;
        RECT 5.465 -0.085 5.715 0.755 ;
        RECT 4.485 -0.085 4.815 0.755 ;
        RECT 3.625 -0.085 3.875 0.755 ;
        RECT 2.845 -0.085 3.015 1.095 ;
        RECT 1.905 -0.085 2.155 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 10.095 2.105 10.425 3.415 ;
        RECT 5.385 2.105 5.555 3.415 ;
        RECT 4.525 2.105 4.695 3.415 ;
        RECT 3.665 2.105 3.835 3.415 ;
        RECT 2.775 2.025 2.945 3.415 ;
        RECT 1.915 2.365 2.085 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.195 0.925 6.225 1.095 ;
      RECT 5.895 0.255 6.225 1.095 ;
      RECT 5.035 0.255 5.285 1.095 ;
      RECT 4.055 0.255 4.305 1.095 ;
      RECT 3.195 0.255 3.445 1.095 ;
      RECT 9.695 0.255 9.945 0.755 ;
      RECT 8.685 0.255 9.015 0.755 ;
      RECT 7.685 0.255 8.015 0.755 ;
      RECT 6.755 0.255 7.085 0.755 ;
      RECT 5.895 0.255 9.945 0.425 ;
      RECT 5.735 2.905 9.915 3.075 ;
      RECT 9.745 2.105 9.915 3.075 ;
      RECT 4.875 1.765 5.205 3.075 ;
      RECT 4.015 1.765 4.345 3.075 ;
      RECT 3.155 1.765 3.485 3.075 ;
      RECT 8.735 2.105 9.065 3.075 ;
      RECT 7.735 2.105 8.065 3.075 ;
      RECT 6.735 2.105 7.065 3.075 ;
      RECT 5.735 1.765 6.065 3.075 ;
      RECT 3.155 1.765 6.065 1.935 ;
      RECT 0.115 1.685 0.365 3.075 ;
      RECT 0.195 0.255 0.365 3.075 ;
      RECT 1.055 1.685 1.225 2.735 ;
      RECT 0.115 1.685 2.985 1.855 ;
      RECT 2.815 1.265 2.985 1.855 ;
      RECT 2.815 1.265 9.82 1.595 ;
      RECT 0.115 0.255 0.365 1.095 ;
      RECT 0.115 0.84 1.375 1.01 ;
      RECT 1.045 0.595 1.375 1.01 ;
      RECT 2.335 0.255 2.665 1.015 ;
      RECT 1.555 0.775 2.665 1.01 ;
      RECT 1.555 0.255 1.725 1.01 ;
      RECT 0.545 0.255 0.875 0.67 ;
      RECT 0.545 0.255 1.725 0.425 ;
      RECT 2.265 2.025 2.595 3.075 ;
      RECT 0.545 2.905 1.735 3.075 ;
      RECT 1.405 2.025 1.735 3.075 ;
      RECT 0.545 2.025 0.875 3.075 ;
      RECT 1.405 2.025 2.595 2.195 ;
  END
END scs130lp_buflp_8

MACRO scs130lp_buflp_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_buflp_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.55 1.795 2.89 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.44 0.475 2.89 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.935 -0.085 1.265 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.965 2.43 1.295 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.965 0.58 2.215 2.89 ;
      RECT 0.66 1.21 0.99 1.88 ;
      RECT 0.66 1.21 2.215 1.38 ;
      RECT 1.755 0.58 2.215 1.38 ;
  END
END scs130lp_buflp_m

MACRO scs130lp_busdriver2_20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busdriver2_20 0 0 ;
  SIZE 24.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.016 LAYER li ;
    PORT
      LAYER li ;
        RECT 21.83 1.18 24.835 1.515 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 1.18 0.445 1.515 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.2502 LAYER li ;
    PORT
      LAYER li ;
        RECT 20.57 1.495 20.82 2.805 ;
        RECT 11.305 1.505 20.82 1.725 ;
        RECT 16.27 1.495 20.82 1.725 ;
        RECT 19.7 1.495 19.89 2.715 ;
        RECT 18.84 1.495 19.03 2.715 ;
        RECT 17.98 1.495 18.17 2.715 ;
        RECT 17.12 1.495 17.31 2.715 ;
        RECT 16.26 1.505 16.45 2.715 ;
        RECT 15.4 1.505 15.59 2.715 ;
        RECT 9.75 0.645 15.4 0.895 ;
        RECT 14.54 1.505 14.73 2.715 ;
        RECT 13.68 1.505 13.87 2.715 ;
        RECT 12.82 1.505 13.01 2.715 ;
        RECT 11.305 1.505 13.01 1.78 ;
        RECT 11.305 0.645 12.235 1.78 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 24.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 24.96 0.085 ;
        RECT 23.56 -0.085 23.89 1 ;
        RECT 22.54 -0.085 22.87 0.65 ;
        RECT 21.52 -0.085 21.85 0.65 ;
        RECT 8.89 -0.085 9.06 0.815 ;
        RECT 8.03 -0.085 8.2 0.815 ;
        RECT 7.17 -0.085 7.34 0.815 ;
        RECT 6.15 -0.085 6.48 0.475 ;
        RECT 5.13 -0.085 5.46 0.475 ;
        RECT 4.27 -0.085 4.6 0.475 ;
        RECT 3.41 -0.085 3.74 0.475 ;
        RECT 2.34 -0.085 2.67 0.445 ;
        RECT 1.055 -0.085 1.385 0.445 ;
        RECT 0.115 -0.085 0.445 1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 24.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 24.96 3.415 ;
        RECT 24.595 1.815 24.845 3.415 ;
        RECT 23.71 2.045 23.88 3.415 ;
        RECT 22.85 2.045 23.02 3.415 ;
        RECT 21.99 2.165 22.16 3.415 ;
        RECT 21.05 1.815 21.3 3.415 ;
        RECT 11.315 2.365 11.645 3.415 ;
        RECT 10.535 1.815 10.705 3.415 ;
        RECT 9.665 2.205 9.855 3.415 ;
        RECT 8.805 2.205 8.995 3.415 ;
        RECT 7.925 2.205 8.115 3.415 ;
        RECT 7.065 2.205 7.255 3.415 ;
        RECT 6.205 2.205 6.395 3.415 ;
        RECT 5.345 2.205 5.535 3.415 ;
        RECT 4.485 2.205 4.675 3.415 ;
        RECT 3.625 2.205 3.815 3.415 ;
        RECT 2.775 1.855 2.945 3.415 ;
        RECT 1.915 2.165 2.085 3.415 ;
        RECT 0.975 1.815 1.225 3.415 ;
        RECT 0.115 1.815 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 24.085 1.695 24.415 3.065 ;
      RECT 23.2 1.695 23.53 3.065 ;
      RECT 22.34 1.695 22.67 3.065 ;
      RECT 21.48 1.695 21.81 3.065 ;
      RECT 21.48 1.695 24.415 1.865 ;
      RECT 21.48 0.83 21.65 3.065 ;
      RECT 12.405 1.075 15.455 1.325 ;
      RECT 12.405 1.075 21.65 1.315 ;
      RECT 15.66 0.985 21.65 1.315 ;
      RECT 23.05 0.265 23.38 1 ;
      RECT 21.48 0.83 23.38 1 ;
      RECT 22.03 0.295 22.36 1 ;
      RECT 12.32 2.885 20.39 3.065 ;
      RECT 20.06 1.895 20.39 3.065 ;
      RECT 10.885 1.465 11.135 3.065 ;
      RECT 10.025 1.465 10.355 3.065 ;
      RECT 19.2 1.895 19.53 3.065 ;
      RECT 18.34 1.895 18.67 3.065 ;
      RECT 17.48 1.895 17.81 3.065 ;
      RECT 16.62 1.895 16.95 3.065 ;
      RECT 15.76 1.895 16.09 3.065 ;
      RECT 14.9 1.895 15.23 3.065 ;
      RECT 14.04 1.895 14.37 3.065 ;
      RECT 13.18 1.895 13.51 3.065 ;
      RECT 12.32 1.96 12.65 3.065 ;
      RECT 9.165 1.865 9.495 2.765 ;
      RECT 8.305 1.865 8.635 2.765 ;
      RECT 7.425 1.865 7.755 2.765 ;
      RECT 6.565 1.865 6.895 2.765 ;
      RECT 5.705 1.865 6.035 2.765 ;
      RECT 4.845 1.865 5.175 2.765 ;
      RECT 3.985 1.865 4.315 2.765 ;
      RECT 3.125 1.865 3.455 2.765 ;
      RECT 10.885 1.96 12.65 2.185 ;
      RECT 3.125 1.865 10.355 2.035 ;
      RECT 10.025 1.465 11.135 1.635 ;
      RECT 6.66 0.995 9.57 1.165 ;
      RECT 9.24 0.265 9.57 1.165 ;
      RECT 8.38 0.265 8.71 1.165 ;
      RECT 7.52 0.265 7.85 1.165 ;
      RECT 6.66 0.265 6.99 1.165 ;
      RECT 2.9 0.655 6.99 0.825 ;
      RECT 15.58 0.265 15.91 0.805 ;
      RECT 5.64 0.265 5.97 0.825 ;
      RECT 4.78 0.265 4.95 0.825 ;
      RECT 3.92 0.265 4.09 0.825 ;
      RECT 2.9 0.265 3.23 0.825 ;
      RECT 9.24 0.265 15.91 0.475 ;
      RECT 2.265 1.515 2.595 3.065 ;
      RECT 1.405 1.815 1.735 3.065 ;
      RECT 1.405 1.815 2.595 1.985 ;
      RECT 1.68 0.975 2.01 1.985 ;
      RECT 2.265 1.515 9.78 1.685 ;
      RECT 6.39 1.345 9.78 1.685 ;
      RECT 0.625 0.265 0.795 3.065 ;
      RECT 2.19 1.005 6.15 1.335 ;
      RECT 2.19 0.625 2.36 1.335 ;
      RECT 0.625 0.625 2.36 0.795 ;
  END
END scs130lp_busdriver2_20

MACRO scs130lp_busdriver_20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busdriver_20 0 0 ;
  SIZE 24.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.016 LAYER li ;
    PORT
      LAYER li ;
        RECT 21.83 1.18 24.835 1.515 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 1.18 0.445 1.515 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.2502 LAYER li ;
    PORT
      LAYER li ;
        RECT 20.57 1.495 20.82 2.805 ;
        RECT 16.27 1.495 20.82 1.665 ;
        RECT 19.71 1.495 19.88 2.715 ;
        RECT 18.85 1.495 19.02 2.715 ;
        RECT 17.99 1.495 18.16 2.715 ;
        RECT 17.13 1.495 17.3 2.715 ;
        RECT 16.27 1.495 16.44 2.715 ;
        RECT 11.305 1.505 16.44 1.675 ;
        RECT 15.41 1.505 15.58 2.715 ;
        RECT 9.75 0.645 15.4 0.895 ;
        RECT 14.55 1.505 14.72 2.715 ;
        RECT 13.69 1.505 13.86 2.715 ;
        RECT 12.83 1.505 13 2.715 ;
        RECT 11.305 1.505 13 1.78 ;
        RECT 11.305 0.645 12.235 1.78 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 24.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 24.96 0.085 ;
        RECT 23.56 -0.085 23.89 1 ;
        RECT 22.54 -0.085 22.87 0.65 ;
        RECT 21.52 -0.085 21.85 0.65 ;
        RECT 8.89 -0.085 9.06 0.815 ;
        RECT 8.03 -0.085 8.2 0.815 ;
        RECT 7.17 -0.085 7.34 0.815 ;
        RECT 6.15 -0.085 6.48 0.475 ;
        RECT 5.13 -0.085 5.46 0.475 ;
        RECT 4.27 -0.085 4.6 0.475 ;
        RECT 3.41 -0.085 3.74 0.475 ;
        RECT 2.34 -0.085 2.67 0.445 ;
        RECT 1.055 -0.085 1.385 0.445 ;
        RECT 0.115 -0.085 0.445 1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 24.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 24.96 3.415 ;
        RECT 24.595 1.815 24.845 3.415 ;
        RECT 23.71 2.045 23.88 3.415 ;
        RECT 22.85 2.045 23.02 3.415 ;
        RECT 21.99 2.165 22.16 3.415 ;
        RECT 21.05 1.815 21.3 3.415 ;
        RECT 11.315 2.365 11.645 3.415 ;
        RECT 10.535 1.815 10.705 3.415 ;
        RECT 9.665 2.205 9.855 3.415 ;
        RECT 8.805 2.205 8.995 3.415 ;
        RECT 7.925 2.205 8.115 3.415 ;
        RECT 7.065 2.205 7.255 3.415 ;
        RECT 6.205 2.205 6.395 3.415 ;
        RECT 5.345 2.205 5.535 3.415 ;
        RECT 4.485 2.205 4.675 3.415 ;
        RECT 3.625 2.205 3.815 3.415 ;
        RECT 2.775 1.855 2.945 3.415 ;
        RECT 1.915 2.165 2.085 3.415 ;
        RECT 0.975 1.815 1.225 3.415 ;
        RECT 0.115 1.815 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 24.085 1.695 24.415 3.065 ;
      RECT 23.2 1.695 23.53 3.065 ;
      RECT 22.34 1.695 22.67 3.065 ;
      RECT 21.48 1.695 21.81 3.065 ;
      RECT 21.48 1.695 24.415 1.865 ;
      RECT 21.48 0.83 21.65 3.065 ;
      RECT 12.405 1.075 15.455 1.325 ;
      RECT 12.405 1.075 21.65 1.315 ;
      RECT 15.66 0.985 21.65 1.315 ;
      RECT 23.05 0.265 23.38 1 ;
      RECT 21.48 0.83 23.38 1 ;
      RECT 22.03 0.295 22.36 1 ;
      RECT 12.32 2.895 20.39 3.065 ;
      RECT 20.06 1.845 20.39 3.065 ;
      RECT 10.885 1.465 11.135 3.065 ;
      RECT 10.025 1.465 10.355 3.065 ;
      RECT 19.2 1.845 19.53 3.065 ;
      RECT 18.34 1.845 18.67 3.065 ;
      RECT 17.48 1.845 17.81 3.065 ;
      RECT 16.62 1.845 16.95 3.065 ;
      RECT 15.76 1.855 16.09 3.065 ;
      RECT 14.9 1.855 15.23 3.065 ;
      RECT 14.04 1.855 14.37 3.065 ;
      RECT 13.18 1.855 13.51 3.065 ;
      RECT 12.32 1.96 12.65 3.065 ;
      RECT 9.165 1.865 9.495 2.765 ;
      RECT 8.305 1.865 8.635 2.765 ;
      RECT 7.425 1.865 7.755 2.765 ;
      RECT 6.565 1.865 6.895 2.765 ;
      RECT 5.705 1.865 6.035 2.765 ;
      RECT 4.845 1.865 5.175 2.765 ;
      RECT 3.985 1.865 4.315 2.765 ;
      RECT 3.125 1.865 3.455 2.765 ;
      RECT 10.885 1.96 12.65 2.185 ;
      RECT 3.125 1.865 10.355 2.035 ;
      RECT 10.025 1.465 11.135 1.635 ;
      RECT 6.66 0.995 9.57 1.165 ;
      RECT 9.24 0.265 9.57 1.165 ;
      RECT 8.38 0.265 8.71 1.165 ;
      RECT 7.52 0.265 7.85 1.165 ;
      RECT 6.66 0.265 6.99 1.165 ;
      RECT 2.9 0.655 6.99 0.825 ;
      RECT 15.58 0.265 15.91 0.805 ;
      RECT 5.64 0.265 5.97 0.825 ;
      RECT 4.78 0.265 4.95 0.825 ;
      RECT 3.92 0.265 4.09 0.825 ;
      RECT 2.9 0.265 3.23 0.825 ;
      RECT 9.24 0.265 15.91 0.475 ;
      RECT 2.265 1.515 2.595 3.065 ;
      RECT 1.405 1.815 1.735 3.065 ;
      RECT 1.405 1.815 2.595 1.985 ;
      RECT 1.68 0.975 2.01 1.985 ;
      RECT 2.265 1.515 9.78 1.685 ;
      RECT 6.39 1.345 9.78 1.685 ;
      RECT 0.625 0.265 0.795 3.065 ;
      RECT 2.19 1.005 6.15 1.335 ;
      RECT 2.19 0.625 2.36 1.335 ;
      RECT 0.625 0.625 2.36 0.795 ;
  END
END scs130lp_busdriver_20

MACRO scs130lp_busdrivernovlp2_20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busdrivernovlp2_20 0 0 ;
  SIZE 17.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.925 1.345 5.255 1.675 ;
        RECT 4.925 1.345 5.155 2.15 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.815 0.995 6.215 1.325 ;
        RECT 5.815 0.645 5.985 1.325 ;
        RECT 4.035 0.645 5.985 0.815 ;
        RECT 4.035 0.265 4.205 0.815 ;
        RECT 3.335 0.265 4.205 0.435 ;
        RECT 2.475 0.85 3.505 1.02 ;
        RECT 3.335 0.265 3.505 1.02 ;
        RECT 2.475 0.265 2.805 1.02 ;
        RECT 1.57 0.265 2.805 0.435 ;
        RECT 0.505 0.995 1.74 1.165 ;
        RECT 1.57 0.265 1.74 1.165 ;
        RECT 0.505 0.995 0.835 1.41 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3528 LAYER li ;
    ANTENNADIFFAREA 4.968 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 9.16 1.92 17.19 2.15 ;
      LAYER li ;
        RECT 16.88 1.94 17.21 3.065 ;
        RECT 16.02 0.255 16.35 3.065 ;
        RECT 15.16 0.26 15.49 3.065 ;
        RECT 14.3 0.255 14.63 3.065 ;
        RECT 13.44 0.255 13.77 3.065 ;
        RECT 12.58 0.255 12.91 3.065 ;
        RECT 11.72 0.255 12.05 3.065 ;
        RECT 10.86 0.255 11.19 3.065 ;
        RECT 10 0.255 10.33 3.065 ;
        RECT 9.22 1.95 10.33 2.13 ;
        RECT 9.22 1.95 9.39 3.065 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 17.76 0.085 ;
        RECT 15.67 -0.085 15.84 0.865 ;
        RECT 14.81 -0.085 14.98 0.865 ;
        RECT 13.95 -0.085 14.12 0.865 ;
        RECT 13.09 -0.085 13.26 0.865 ;
        RECT 12.23 -0.085 12.4 0.865 ;
        RECT 11.37 -0.085 11.54 0.865 ;
        RECT 10.51 -0.085 10.68 0.865 ;
        RECT 7.745 -0.085 7.995 0.745 ;
        RECT 6.675 -0.085 7.005 0.465 ;
        RECT 5.545 -0.085 5.875 0.465 ;
        RECT 4.385 -0.085 4.715 0.465 ;
        RECT 2.985 -0.085 3.155 0.67 ;
        RECT 1.06 -0.085 1.39 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 17.76 3.415 ;
        RECT 17.39 2.29 17.64 3.415 ;
        RECT 16.53 2.29 16.7 3.415 ;
        RECT 15.67 2.29 15.84 3.415 ;
        RECT 14.81 2.29 14.98 3.415 ;
        RECT 13.95 2.29 14.12 3.415 ;
        RECT 13.09 2.29 13.26 3.415 ;
        RECT 12.23 2.29 12.4 3.415 ;
        RECT 11.37 2.29 11.54 3.415 ;
        RECT 10.51 2.29 10.68 3.415 ;
        RECT 9.57 2.31 9.82 3.415 ;
        RECT 8.205 2.135 8.875 3.415 ;
        RECT 7.265 2.185 7.515 3.415 ;
        RECT 5.845 1.845 6.175 3.415 ;
        RECT 4.665 2.68 4.995 3.415 ;
        RECT 2.51 2.435 2.76 3.415 ;
        RECT 1.57 2.29 1.82 3.415 ;
        RECT 0.63 1.94 0.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 9.215 1.55 17.11 1.78 ;
      RECT 2.015 1.55 2.305 1.78 ;
      RECT 2.015 1.595 17.11 1.735 ;
      RECT 9.6 1.18 13.33 1.41 ;
      RECT 6.335 1.18 6.625 1.41 ;
      RECT 5.375 1.18 5.665 1.41 ;
      RECT 5.375 1.225 13.33 1.365 ;
    LAYER li ;
      RECT 7.695 1.785 8.025 3.065 ;
      RECT 7.695 1.785 9.04 1.955 ;
      RECT 8.87 0.615 9.04 1.955 ;
      RECT 8.87 1.55 9.475 1.78 ;
      RECT 8.685 0.615 9.04 1.095 ;
      RECT 9.22 0.265 9.47 1.095 ;
      RECT 7.36 0.925 8.505 1.095 ;
      RECT 8.175 0.265 8.505 1.095 ;
      RECT 7.36 0.295 7.565 1.095 ;
      RECT 7.235 0.295 7.565 0.465 ;
      RECT 8.175 0.265 9.47 0.435 ;
      RECT 6.665 1.845 6.995 2.725 ;
      RECT 6.665 1.845 7.19 2.015 ;
      RECT 7.02 0.645 7.19 2.015 ;
      RECT 7.02 1.275 8.69 1.605 ;
      RECT 6.165 0.645 7.19 0.815 ;
      RECT 6.165 0.265 6.495 0.815 ;
      RECT 3.685 1.815 3.975 2.715 ;
      RECT 3.685 0.615 3.855 2.715 ;
      RECT 5.435 0.995 5.635 1.41 ;
      RECT 3.685 0.995 5.635 1.165 ;
      RECT 5.335 1.855 5.585 3.065 ;
      RECT 3.335 2.895 4.485 3.065 ;
      RECT 4.155 1.815 4.485 3.065 ;
      RECT 3.335 1.815 3.505 3.065 ;
      RECT 4.155 2.33 5.585 2.5 ;
      RECT 2 2.085 2.33 3.065 ;
      RECT 2 2.085 3.13 2.255 ;
      RECT 2.8 1.575 3.13 2.255 ;
      RECT 2.8 1.2 2.97 2.255 ;
      RECT 1.995 1.2 2.97 1.37 ;
      RECT 1.995 0.615 2.245 1.37 ;
      RECT 1.06 1.94 1.39 3.065 ;
      RECT 1.06 1.94 1.765 2.11 ;
      RECT 1.595 1.55 1.765 2.11 ;
      RECT 2.045 1.55 2.565 1.905 ;
      RECT 1.595 1.55 2.565 1.72 ;
      RECT 0.1 1.59 0.43 2.695 ;
      RECT 0.1 1.59 1.415 1.76 ;
      RECT 1.085 1.345 1.415 1.76 ;
      RECT 0.1 0.645 0.27 2.695 ;
      RECT 0.1 0.645 0.88 0.815 ;
      RECT 0.55 0.405 0.88 0.815 ;
      RECT 16.52 1.345 17.11 1.76 ;
      RECT 15.66 1.345 15.85 1.76 ;
      RECT 14.8 1.345 14.99 1.76 ;
      RECT 13.94 1.345 14.13 1.76 ;
      RECT 13.08 1.035 13.27 1.41 ;
      RECT 12.22 1.035 12.41 1.41 ;
      RECT 11.36 1.035 11.55 1.41 ;
      RECT 10.5 1.035 10.69 1.41 ;
      RECT 9.64 1.035 9.83 1.41 ;
      RECT 6.395 0.995 6.84 1.665 ;
  END
END scs130lp_busdrivernovlp2_20

MACRO scs130lp_busdrivernovlp_20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busdrivernovlp_20 0 0 ;
  SIZE 17.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.925 1.345 5.255 1.675 ;
        RECT 4.925 1.345 5.155 2.15 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.815 0.995 6.215 1.325 ;
        RECT 5.815 0.645 5.985 1.325 ;
        RECT 4.035 0.645 5.985 0.815 ;
        RECT 4.035 0.265 4.205 0.815 ;
        RECT 3.335 0.265 4.205 0.435 ;
        RECT 2.475 0.85 3.505 1.02 ;
        RECT 3.335 0.265 3.505 1.02 ;
        RECT 2.475 0.265 2.805 1.02 ;
        RECT 1.57 0.265 2.805 0.435 ;
        RECT 0.505 0.995 1.74 1.165 ;
        RECT 1.57 0.265 1.74 1.165 ;
        RECT 0.505 0.995 0.835 1.41 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3528 LAYER li ;
    ANTENNADIFFAREA 4.968 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 9.16 1.92 17.19 2.15 ;
      LAYER li ;
        RECT 16.88 1.94 17.21 3.065 ;
        RECT 16.02 0.255 16.35 3.065 ;
        RECT 15.16 0.26 15.49 3.065 ;
        RECT 14.3 0.255 14.63 3.065 ;
        RECT 13.44 0.255 13.77 3.065 ;
        RECT 12.58 0.255 12.91 3.065 ;
        RECT 11.72 0.255 12.05 3.065 ;
        RECT 10.86 0.255 11.19 3.065 ;
        RECT 10 0.255 10.33 3.065 ;
        RECT 9.22 1.95 10.33 2.13 ;
        RECT 9.22 1.95 9.39 3.065 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 17.76 0.085 ;
        RECT 15.67 -0.085 15.84 0.865 ;
        RECT 14.81 -0.085 14.98 0.865 ;
        RECT 13.95 -0.085 14.12 0.865 ;
        RECT 13.09 -0.085 13.26 0.865 ;
        RECT 12.23 -0.085 12.4 0.865 ;
        RECT 11.37 -0.085 11.54 0.865 ;
        RECT 10.51 -0.085 10.68 0.865 ;
        RECT 7.745 -0.085 7.995 0.745 ;
        RECT 6.675 -0.085 7.005 0.465 ;
        RECT 5.545 -0.085 5.875 0.465 ;
        RECT 4.385 -0.085 4.715 0.465 ;
        RECT 2.985 -0.085 3.155 0.67 ;
        RECT 1.06 -0.085 1.39 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 17.76 3.415 ;
        RECT 17.39 2.29 17.64 3.415 ;
        RECT 16.53 2.29 16.7 3.415 ;
        RECT 15.67 2.29 15.84 3.415 ;
        RECT 14.81 2.29 14.98 3.415 ;
        RECT 13.95 2.29 14.12 3.415 ;
        RECT 13.09 2.29 13.26 3.415 ;
        RECT 12.23 2.29 12.4 3.415 ;
        RECT 11.37 2.29 11.54 3.415 ;
        RECT 10.51 2.29 10.68 3.415 ;
        RECT 9.57 2.31 9.82 3.415 ;
        RECT 8.205 2.135 8.875 3.415 ;
        RECT 7.265 2.185 7.515 3.415 ;
        RECT 5.845 1.845 6.175 3.415 ;
        RECT 4.665 2.68 4.995 3.415 ;
        RECT 2.51 2.435 2.76 3.415 ;
        RECT 1.57 2.29 1.82 3.415 ;
        RECT 0.63 1.94 0.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 9.215 1.55 17.11 1.78 ;
      RECT 2.015 1.55 2.305 1.78 ;
      RECT 2.015 1.595 17.11 1.735 ;
      RECT 9.6 1.18 13.33 1.41 ;
      RECT 6.335 1.18 6.625 1.41 ;
      RECT 5.375 1.18 5.665 1.41 ;
      RECT 5.375 1.225 13.33 1.365 ;
    LAYER li ;
      RECT 7.695 1.785 8.025 3.065 ;
      RECT 7.695 1.785 9.04 1.955 ;
      RECT 8.87 0.615 9.04 1.955 ;
      RECT 8.87 1.55 9.475 1.78 ;
      RECT 8.685 0.615 9.04 1.095 ;
      RECT 9.22 0.265 9.47 1.095 ;
      RECT 7.36 0.925 8.505 1.095 ;
      RECT 8.175 0.265 8.505 1.095 ;
      RECT 7.36 0.295 7.565 1.095 ;
      RECT 7.235 0.295 7.565 0.465 ;
      RECT 8.175 0.265 9.47 0.435 ;
      RECT 6.665 1.845 6.995 2.725 ;
      RECT 6.665 1.845 7.19 2.015 ;
      RECT 7.02 0.645 7.19 2.015 ;
      RECT 7.02 1.275 8.69 1.605 ;
      RECT 6.165 0.645 7.19 0.815 ;
      RECT 6.165 0.265 6.495 0.815 ;
      RECT 3.685 1.815 3.975 2.715 ;
      RECT 3.685 0.615 3.855 2.715 ;
      RECT 5.435 0.995 5.635 1.41 ;
      RECT 3.685 0.995 5.635 1.165 ;
      RECT 5.335 1.855 5.585 3.065 ;
      RECT 3.335 2.895 4.485 3.065 ;
      RECT 4.155 1.815 4.485 3.065 ;
      RECT 3.335 1.815 3.505 3.065 ;
      RECT 4.155 2.33 5.585 2.5 ;
      RECT 2 2.085 2.33 3.065 ;
      RECT 2 2.085 3.13 2.255 ;
      RECT 2.8 1.575 3.13 2.255 ;
      RECT 2.8 1.2 2.97 2.255 ;
      RECT 1.995 1.2 2.97 1.37 ;
      RECT 1.995 0.615 2.245 1.37 ;
      RECT 1.06 1.94 1.39 3.065 ;
      RECT 1.06 1.94 1.765 2.11 ;
      RECT 1.595 1.55 1.765 2.11 ;
      RECT 2.045 1.55 2.565 1.905 ;
      RECT 1.595 1.55 2.565 1.72 ;
      RECT 0.1 1.59 0.43 2.695 ;
      RECT 0.1 1.59 1.415 1.76 ;
      RECT 1.085 1.345 1.415 1.76 ;
      RECT 0.1 0.645 0.27 2.695 ;
      RECT 0.1 0.645 0.88 0.815 ;
      RECT 0.55 0.405 0.88 0.815 ;
      RECT 16.52 1.345 17.11 1.76 ;
      RECT 15.66 1.345 15.85 1.76 ;
      RECT 14.8 1.345 14.99 1.76 ;
      RECT 13.94 1.345 14.13 1.76 ;
      RECT 13.08 1.035 13.27 1.41 ;
      RECT 12.22 1.035 12.41 1.41 ;
      RECT 11.36 1.035 11.55 1.41 ;
      RECT 10.5 1.035 10.69 1.41 ;
      RECT 9.64 1.035 9.83 1.41 ;
      RECT 6.395 0.995 6.84 1.665 ;
  END
END scs130lp_busdrivernovlp_20

MACRO scs130lp_busdrivernovlpsleep_20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busdrivernovlpsleep_20 0 0 ;
  SIZE 23.52 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.4 0.44 12.385 0.77 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.348 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.2 2.415 1.59 ;
    END
  END TEB
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 1.228 LAYER met1 ;
      ANTENNAMAXAREACAR 1.253571 LAYER li ;
      ANTENNAMAXAREACAR 1.253571 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.261905 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.261905 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 11.72 1.92 12.01 2.15 ;
        RECT 0.625 1.95 12.01 2.12 ;
        RECT 5.355 1.92 5.645 2.15 ;
        RECT 0.625 1.92 0.915 2.15 ;
      LAYER li ;
        RECT 11.445 1.325 12.115 1.615 ;
        RECT 11.71 1.325 12.055 2.15 ;
        RECT 5.27 1.765 5.675 2.155 ;
        RECT 0.595 1.2 0.925 2.15 ;
    END
  END SLEEP
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3528 LAYER li ;
    ANTENNADIFFAREA 4.968 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 14.48 1.92 22.51 2.15 ;
      LAYER li ;
        RECT 22.2 1.94 22.53 3.065 ;
        RECT 21.34 0.255 21.67 3.065 ;
        RECT 20.48 0.26 20.81 3.065 ;
        RECT 19.62 0.255 19.95 3.065 ;
        RECT 18.76 0.255 19.09 3.065 ;
        RECT 17.9 0.255 18.23 3.065 ;
        RECT 17.04 0.255 17.37 3.065 ;
        RECT 16.18 0.255 16.51 3.065 ;
        RECT 15.32 0.255 15.65 3.065 ;
        RECT 14.54 1.95 15.65 2.13 ;
        RECT 14.54 1.95 14.71 3.065 ;
    END
  END Z
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 23.45 2.945 ;
      LAYER li ;
        RECT 4.885 2.665 5.215 3.015 ;
        RECT 4.065 1.85 4.315 3.045 ;
        RECT 2.495 2.44 3.4 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 23.52 0.245 ;
      LAYER li ;
        RECT 0 -0.085 23.52 0.085 ;
        RECT 20.99 -0.085 21.16 0.865 ;
        RECT 20.13 -0.085 20.3 0.865 ;
        RECT 19.27 -0.085 19.44 0.865 ;
        RECT 18.41 -0.085 18.58 0.865 ;
        RECT 17.55 -0.085 17.72 0.865 ;
        RECT 16.69 -0.085 16.86 0.865 ;
        RECT 15.83 -0.085 16 0.865 ;
        RECT 13.055 -0.085 13.365 0.755 ;
        RECT 10.72 -0.085 11.05 0.465 ;
        RECT 9.455 -0.085 10.19 0.485 ;
        RECT 8.415 -0.085 8.785 0.465 ;
        RECT 6.975 -0.085 7.225 0.68 ;
        RECT 3.675 -0.085 5.11 0.475 ;
        RECT 2.72 -0.085 2.995 1.04 ;
        RECT 1.805 -0.085 2.135 0.69 ;
        RECT 0.945 -0.085 1.25 1.02 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 23.52 3.575 ;
      LAYER li ;
        RECT 0 3.245 23.52 3.415 ;
        RECT 22.71 2.29 22.96 3.415 ;
        RECT 21.85 2.29 22.02 3.415 ;
        RECT 20.99 2.29 21.16 3.415 ;
        RECT 20.13 2.29 20.3 3.415 ;
        RECT 19.27 2.29 19.44 3.415 ;
        RECT 18.41 2.29 18.58 3.415 ;
        RECT 17.55 2.29 17.72 3.415 ;
        RECT 16.69 2.29 16.86 3.415 ;
        RECT 15.83 2.29 16 3.415 ;
        RECT 14.89 2.31 15.14 3.415 ;
        RECT 14.025 2.135 14.36 3.415 ;
        RECT 12.2 2.735 12.46 3.415 ;
        RECT 11.27 2.32 11.53 3.415 ;
        RECT 9.71 1.845 10.04 3.415 ;
        RECT 8.78 2.67 9.04 3.415 ;
        RECT 6.705 2.435 6.955 3.415 ;
        RECT 5.405 2.665 5.735 3.415 ;
        RECT 0.625 2.32 0.955 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 14.5 1.595 22.465 1.78 ;
      RECT 14.505 1.55 22.465 1.78 ;
      RECT 6.335 1.55 6.625 1.78 ;
      RECT 6.335 1.595 22.465 1.735 ;
      RECT 14.92 1.18 18.695 1.41 ;
      RECT 10.425 1.18 10.715 1.41 ;
      RECT 9.455 1.18 9.745 1.41 ;
      RECT 9.455 1.225 18.695 1.365 ;
      RECT 4.505 1.55 4.795 1.78 ;
      RECT 0.095 1.55 0.385 1.78 ;
      RECT 0.095 1.595 4.795 1.735 ;
    LAYER li ;
      RECT 13.15 1.785 13.41 2.605 ;
      RECT 13.15 1.785 14.37 1.955 ;
      RECT 14.2 0.615 14.37 1.955 ;
      RECT 14.2 1.55 14.86 1.78 ;
      RECT 14.075 0.615 14.37 1.095 ;
      RECT 14.54 0.265 14.79 1.095 ;
      RECT 12.68 0.925 13.905 1.095 ;
      RECT 13.575 0.265 13.905 1.095 ;
      RECT 12.68 0.295 12.885 1.095 ;
      RECT 12.555 0.295 12.885 0.465 ;
      RECT 13.575 0.265 14.79 0.435 ;
      RECT 10.5 1.845 10.83 2.725 ;
      RECT 10.5 1.845 11.14 2.015 ;
      RECT 10.97 0.645 11.14 2.015 ;
      RECT 12.285 1.275 14.03 1.605 ;
      RECT 12.285 0.955 12.455 1.605 ;
      RECT 10.97 0.955 12.455 1.13 ;
      RECT 10.36 0.645 11.14 0.815 ;
      RECT 10.36 0.265 10.55 0.815 ;
      RECT 12.65 2.775 13.84 3.075 ;
      RECT 13.59 2.185 13.84 3.075 ;
      RECT 11.7 2.32 12.03 3.035 ;
      RECT 12.65 2.185 12.98 3.075 ;
      RECT 11.7 2.32 12.98 2.49 ;
      RECT 1.995 2.1 2.325 3.075 ;
      RECT 1.995 2.1 3.505 2.27 ;
      RECT 3.335 0.275 3.505 2.27 ;
      RECT 9.985 0.995 10.315 1.325 ;
      RECT 6.525 0.85 7.565 1.02 ;
      RECT 7.395 0.265 7.565 1.02 ;
      RECT 9.985 0.655 10.155 1.325 ;
      RECT 6.525 0.265 6.695 1.02 ;
      RECT 8.075 0.655 10.155 0.825 ;
      RECT 3.335 0.645 5.455 0.815 ;
      RECT 5.285 0.265 5.455 0.815 ;
      RECT 8.075 0.265 8.245 0.825 ;
      RECT 3.185 0.275 3.505 0.605 ;
      RECT 7.395 0.265 8.245 0.435 ;
      RECT 5.285 0.265 6.695 0.435 ;
      RECT 7.92 0.995 8.11 2.715 ;
      RECT 9.455 0.995 9.745 1.505 ;
      RECT 7.735 0.995 8.11 1.225 ;
      RECT 7.735 0.995 9.745 1.165 ;
      RECT 7.735 0.605 7.905 1.225 ;
      RECT 9.21 2.32 9.47 3.065 ;
      RECT 7.5 2.895 8.61 3.065 ;
      RECT 8.28 1.815 8.61 3.065 ;
      RECT 7.5 1.815 7.75 3.065 ;
      RECT 8.28 2.32 9.47 2.5 ;
      RECT 4.485 2.06 4.715 3.07 ;
      RECT 6.195 2.085 6.525 3.065 ;
      RECT 4.485 2.325 6.525 2.495 ;
      RECT 6.195 2.085 7.23 2.255 ;
      RECT 6.97 1.2 7.23 2.255 ;
      RECT 6.185 1.2 7.23 1.37 ;
      RECT 6.185 0.605 6.355 1.37 ;
      RECT 5.66 0.605 6.355 0.815 ;
      RECT 3.675 0.985 3.895 3.065 ;
      RECT 6.335 1.55 6.76 1.905 ;
      RECT 5.845 1.55 6.76 1.72 ;
      RECT 5.845 0.985 6.015 1.72 ;
      RECT 3.675 0.985 6.015 1.155 ;
      RECT 1.475 1.76 1.805 3.065 ;
      RECT 1.42 1.76 3.165 1.93 ;
      RECT 2.9 1.345 3.165 1.93 ;
      RECT 1.42 0.255 1.625 1.93 ;
      RECT 1.42 0.86 2.55 1.03 ;
      RECT 2.305 0.255 2.55 1.03 ;
      RECT 1.42 0.255 1.635 1.03 ;
      RECT 21.84 1.345 22.43 1.76 ;
      RECT 20.98 1.345 21.17 1.76 ;
      RECT 20.12 1.345 20.31 1.76 ;
      RECT 19.26 1.345 19.45 1.76 ;
      RECT 18.4 1.035 18.59 1.41 ;
      RECT 17.54 1.035 17.73 1.41 ;
      RECT 16.68 1.035 16.87 1.41 ;
      RECT 15.82 1.035 16.01 1.41 ;
      RECT 14.96 1.035 15.15 1.41 ;
      RECT 10.485 0.995 10.8 1.665 ;
      RECT 4.485 1.325 4.815 1.815 ;
      RECT 0.095 0.255 0.425 3.075 ;
  END
END scs130lp_busdrivernovlpsleep_20

MACRO scs130lp_bushold0_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bushold0_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.525 1.355 2.195 ;
    END
  END RESET
  PIN X
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 0.84 2.315 3.05 ;
        RECT 0.485 2.365 2.315 2.535 ;
        RECT 1.225 0.84 2.315 1.015 ;
        RECT 1.225 0.255 1.525 1.015 ;
        RECT 0.485 1.525 0.815 2.535 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.975 -0.085 2.305 0.61 ;
        RECT 0.795 -0.085 1.055 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.835 2.72 1.165 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 2.72 0.425 3.05 ;
      RECT 0.085 1.055 0.315 3.05 ;
      RECT 1.605 1.185 1.855 2.195 ;
      RECT 0.085 1.185 1.855 1.355 ;
      RECT 0.085 1.055 0.625 1.355 ;
      RECT 0.335 0.255 0.625 1.355 ;
  END
END scs130lp_bushold0_1

MACRO scs130lp_bushold_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_bushold_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.135 1.355 2.195 ;
    END
  END RESET
  PIN X
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 0.255 2.315 3.05 ;
        RECT 0.485 2.365 2.315 2.535 ;
        RECT 0.485 1.135 0.815 2.535 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.225 -0.085 1.525 0.545 ;
        RECT 0.335 -0.085 0.625 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.195 2.72 1.525 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 2.72 0.735 3.05 ;
      RECT 0.085 0.715 0.315 3.05 ;
      RECT 1.605 0.715 1.855 2.195 ;
      RECT 0.085 0.715 1.855 0.965 ;
      RECT 0.795 0.265 1.055 0.965 ;
  END
END scs130lp_bushold_1

MACRO scs130lp_busreceiver_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busreceiver_0 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.89 1.15 1.345 1.885 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 2.395 0.4 3.075 ;
        RECT 0.09 0.285 0.39 0.615 ;
        RECT 0.09 1.605 0.34 3.075 ;
        RECT 0.09 0.285 0.26 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.56 -0.085 0.89 0.615 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.57 2.395 0.825 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.995 2.055 1.345 3.075 ;
      RECT 0.51 2.055 1.345 2.225 ;
      RECT 0.51 0.785 0.68 2.225 ;
      RECT 0.43 0.785 0.68 1.455 ;
      RECT 0.43 0.785 1.345 0.97 ;
      RECT 1.06 0.3 1.345 0.97 ;
  END
END scs130lp_busreceiver_0

MACRO scs130lp_busreceiver_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busreceiver_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 1.19 1.355 1.435 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.865 0.355 3.075 ;
        RECT 0.085 0.255 0.355 1.03 ;
        RECT 0.085 0.255 0.26 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.525 -0.085 0.855 0.68 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.525 1.945 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.025 1.605 1.345 2.485 ;
      RECT 0.505 1.605 1.345 1.775 ;
      RECT 0.43 1.185 0.695 1.705 ;
      RECT 0.525 0.85 0.695 1.775 ;
      RECT 0.525 0.85 1.345 1.02 ;
      RECT 1.025 0.69 1.345 1.02 ;
  END
END scs130lp_busreceiver_1

MACRO scs130lp_busreceiver_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_busreceiver_m 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 0.875 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.46 0.365 2.96 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.585 -0.085 0.795 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.585 2.76 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.015 1.93 1.225 2.96 ;
      RECT 1.055 0.33 1.225 2.96 ;
      RECT 0.545 1.93 1.225 2.1 ;
      RECT 1.015 0.33 1.225 0.66 ;
  END
END scs130lp_busreceiver_m

MACRO scs130lp_clkbuf_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuf_0 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.89 1.15 1.345 1.885 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 2.395 0.4 3.075 ;
        RECT 0.09 0.285 0.39 0.615 ;
        RECT 0.09 1.605 0.34 3.075 ;
        RECT 0.09 0.285 0.26 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.56 -0.085 0.89 0.615 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.57 2.395 0.825 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.995 2.055 1.285 3.075 ;
      RECT 0.51 2.055 1.285 2.225 ;
      RECT 0.51 0.785 0.68 2.225 ;
      RECT 0.43 0.785 0.68 1.455 ;
      RECT 0.43 0.785 1.345 0.97 ;
      RECT 1.06 0.3 1.345 0.97 ;
  END
END scs130lp_clkbuf_0

MACRO scs130lp_clkbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuf_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.345 1.015 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.3 0.43 0.635 ;
        RECT 0.085 1.525 0.395 3.075 ;
        RECT 0.085 0.3 0.255 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.6 -0.085 0.875 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.565 1.92 0.825 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.995 1.92 1.355 3.075 ;
      RECT 1.185 0.3 1.355 3.075 ;
      RECT 0.425 0.805 1.355 1.135 ;
      RECT 1.045 0.3 1.355 1.135 ;
  END
END scs130lp_clkbuf_1

MACRO scs130lp_clkbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuf_16 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.008 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.43 1.125 1.815 1.455 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    ANTENNADIFFAREA 3.7632 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 2.685 1.92 9.035 2.15 ;
      LAYER li ;
        RECT 8.745 0.275 8.955 3.055 ;
        RECT 7.885 0.275 8.095 3.055 ;
        RECT 7.02 0.275 7.235 3.055 ;
        RECT 6.165 0.275 6.375 3.055 ;
        RECT 5.305 0.275 5.515 3.055 ;
        RECT 4.445 0.275 4.655 3.055 ;
        RECT 3.585 0.275 3.795 3.055 ;
        RECT 2.72 0.275 2.935 3.055 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 9.125 -0.085 9.445 0.605 ;
        RECT 8.265 -0.085 8.575 0.605 ;
        RECT 7.405 -0.085 7.715 0.605 ;
        RECT 6.545 -0.085 6.85 0.605 ;
        RECT 5.685 -0.085 5.995 0.605 ;
        RECT 4.825 -0.085 5.135 0.605 ;
        RECT 3.965 -0.085 4.275 0.605 ;
        RECT 3.105 -0.085 3.415 0.605 ;
        RECT 1.875 -0.085 2.55 0.605 ;
        RECT 1.01 -0.085 1.29 0.605 ;
        RECT 0.125 -0.085 0.42 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 9.125 1.875 9.445 3.415 ;
        RECT 8.265 1.875 8.575 3.415 ;
        RECT 7.405 1.875 7.715 3.415 ;
        RECT 6.545 1.875 6.85 3.415 ;
        RECT 5.685 1.875 5.995 3.415 ;
        RECT 4.825 1.875 5.135 3.415 ;
        RECT 3.965 1.875 4.275 3.415 ;
        RECT 3.105 1.875 3.415 3.415 ;
        RECT 1.88 2.025 2.55 3.415 ;
        RECT 1.025 2.025 1.29 3.415 ;
        RECT 0.125 1.875 0.42 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.96 1.18 8.61 1.41 ;
    LAYER li ;
      RECT 1.46 1.685 1.71 3.075 ;
      RECT 0.59 1.685 0.855 3.075 ;
      RECT 0.59 1.685 2.2 1.855 ;
      RECT 1.985 0.775 2.2 1.855 ;
      RECT 1.985 0.775 2.55 1.535 ;
      RECT 0.59 0.775 2.55 0.945 ;
      RECT 1.46 0.28 1.705 0.945 ;
      RECT 0.59 0.28 0.84 0.945 ;
      RECT 8.265 1.205 8.575 1.535 ;
      RECT 7.405 1.205 7.715 1.535 ;
      RECT 6.545 1.205 6.85 1.535 ;
      RECT 5.685 1.205 5.995 1.535 ;
      RECT 4.825 1.205 5.135 1.535 ;
      RECT 3.965 1.205 4.275 1.535 ;
      RECT 3.105 1.205 3.415 1.535 ;
  END
END scs130lp_clkbuf_16

MACRO scs130lp_clkbuf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuf_2 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.425 0.775 0.875 1.105 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.725 1.815 1.895 ;
        RECT 1.385 0.78 1.815 1.895 ;
        RECT 1.045 0.78 1.815 1.105 ;
        RECT 1.045 1.725 1.305 3.045 ;
        RECT 1.045 0.265 1.305 1.105 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.475 -0.085 1.73 0.61 ;
        RECT 0.555 -0.085 0.83 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.475 2.065 1.73 3.415 ;
        RECT 0.565 1.875 0.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.275 0.395 3.045 ;
      RECT 0.085 1.275 1.215 1.535 ;
      RECT 0.085 0.265 0.255 3.045 ;
      RECT 0.085 0.265 0.385 0.605 ;
  END
END scs130lp_clkbuf_2

MACRO scs130lp_clkbuf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuf_4 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.425 0.775 0.805 1.105 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9408 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.725 2.765 1.895 ;
        RECT 2.255 0.775 2.765 1.895 ;
        RECT 1.045 0.775 2.765 1.025 ;
        RECT 1.905 1.725 2.165 3.06 ;
        RECT 1.905 0.275 2.165 1.025 ;
        RECT 1.045 1.725 1.305 3.06 ;
        RECT 1.045 0.275 1.305 1.025 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.335 -0.085 2.615 0.605 ;
        RECT 1.475 -0.085 1.73 0.605 ;
        RECT 0.555 -0.085 0.83 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.335 2.065 2.62 3.415 ;
        RECT 1.475 2.065 1.73 3.415 ;
        RECT 0.565 1.875 0.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.275 0.395 3.06 ;
      RECT 0.085 1.275 2.085 1.535 ;
      RECT 1.075 1.205 2.085 1.535 ;
      RECT 0.085 0.275 0.255 3.06 ;
      RECT 0.085 0.275 0.385 0.605 ;
  END
END scs130lp_clkbuf_4

MACRO scs130lp_clkbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuf_8 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.4 1.57 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8816 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.42 1.655 4.73 1.895 ;
        RECT 3.76 0.735 4.73 1.895 ;
        RECT 4 0.28 4.26 3.075 ;
        RECT 1.42 0.735 4.73 0.975 ;
        RECT 3.14 1.655 3.4 3.075 ;
        RECT 3.14 0.28 3.4 0.975 ;
        RECT 2.28 1.655 2.54 3.075 ;
        RECT 2.28 0.28 2.54 0.975 ;
        RECT 1.42 1.655 1.68 3.075 ;
        RECT 1.42 0.28 1.68 0.975 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.43 -0.085 4.73 0.565 ;
        RECT 3.57 -0.085 3.83 0.565 ;
        RECT 2.71 -0.085 2.97 0.565 ;
        RECT 1.85 -0.085 2.11 0.565 ;
        RECT 0.99 -0.085 1.25 0.61 ;
        RECT 0.145 -0.085 0.39 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.43 2.065 4.725 3.415 ;
        RECT 3.57 2.065 3.83 3.415 ;
        RECT 2.71 2.065 2.97 3.415 ;
        RECT 1.85 2.065 2.11 3.415 ;
        RECT 0.99 1.875 1.25 3.415 ;
        RECT 0.095 1.875 0.39 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.57 0.265 0.82 3.075 ;
      RECT 0.57 1.155 3.59 1.485 ;
  END
END scs130lp_clkbuf_8

MACRO scs130lp_clkbuf_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuf_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 0.44 1.795 1.485 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.23 1.835 0.56 3.055 ;
        RECT 0.125 0.265 0.495 2.89 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.955 -0.085 1.285 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.76 2.015 1.09 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.535 1.665 1.865 3.055 ;
      RECT 0.74 1.665 2.225 1.835 ;
      RECT 1.975 0.265 2.225 1.835 ;
      RECT 0.74 1.165 1.07 1.835 ;
  END
END scs130lp_clkbuf_lp

MACRO scs130lp_clkbuflp_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuflp_16 0 0 ;
  SIZE 12.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.16 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.775 0.695 1.565 ;
        RECT 0.125 0.775 0.37 1.805 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.28 LAYER li ;
    ANTENNADIFFAREA 3.01 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 3.805 1.92 11.555 2.15 ;
      LAYER li ;
        RECT 11.225 1.92 11.555 3.075 ;
        RECT 10.385 0.265 10.715 1.79 ;
        RECT 10.165 1.17 10.495 3.075 ;
        RECT 9.105 1.17 9.435 3.075 ;
        RECT 8.805 0.265 9.135 1.79 ;
        RECT 8.045 1.92 8.375 3.075 ;
        RECT 7.225 0.265 7.555 1.79 ;
        RECT 6.985 1.17 7.315 3.075 ;
        RECT 5.925 1.17 6.255 3.075 ;
        RECT 5.645 0.265 5.975 1.79 ;
        RECT 4.865 1.92 5.195 3.075 ;
        RECT 4.08 0.265 4.395 1.875 ;
        RECT 3.805 1.705 4.135 3.075 ;
        RECT 4.065 0.265 4.395 1.035 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.48 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.48 0.085 ;
        RECT 11.175 -0.085 11.505 0.605 ;
        RECT 9.595 -0.085 9.925 0.605 ;
        RECT 8.015 -0.085 8.345 0.605 ;
        RECT 6.435 -0.085 6.765 0.605 ;
        RECT 4.855 -0.085 5.185 0.605 ;
        RECT 3.255 -0.085 3.585 0.605 ;
        RECT 1.675 -0.085 2.005 0.605 ;
        RECT 0.125 -0.085 0.425 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.48 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.48 3.415 ;
        RECT 11.755 2.085 12.085 3.415 ;
        RECT 10.695 2.085 11.025 3.415 ;
        RECT 9.635 2.085 9.965 3.415 ;
        RECT 8.575 2.085 8.905 3.415 ;
        RECT 7.515 2.085 7.845 3.415 ;
        RECT 6.455 2.085 6.785 3.415 ;
        RECT 5.395 2.085 5.725 3.415 ;
        RECT 4.335 2.085 4.665 3.415 ;
        RECT 3.275 2.085 3.605 3.415 ;
        RECT 2.215 2.085 2.545 3.415 ;
        RECT 1.225 2.065 1.485 3.415 ;
        RECT 0.095 2.065 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 2.975 1.18 11.905 1.41 ;
    LAYER li ;
      RECT 2.745 1.18 3.075 3.075 ;
      RECT 1.685 1.205 2.015 3.075 ;
      RECT 0.595 2.015 1.055 3.075 ;
      RECT 0.885 0.265 1.055 3.075 ;
      RECT 0.885 1.205 3.91 1.535 ;
      RECT 2.45 1.18 3.91 1.535 ;
      RECT 0.885 0.265 1.23 1.535 ;
      RECT 2.45 0.265 2.795 1.535 ;
      RECT 10.91 1.18 11.92 1.51 ;
      RECT 9.65 1.18 9.98 1.51 ;
      RECT 7.75 1.18 8.555 1.51 ;
      RECT 6.47 1.18 6.8 1.51 ;
      RECT 4.585 1.18 5.39 1.51 ;
  END
END scs130lp_clkbuflp_16

MACRO scs130lp_clkbuflp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuflp_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 0.775 1.325 1.105 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3976 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.555 0.265 2.27 1.875 ;
        RECT 1.32 1.705 1.68 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.465 -0.085 2.795 0.605 ;
        RECT 0.885 -0.085 1.215 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.88 2.085 2.21 3.415 ;
        RECT 0.82 2.065 1.15 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.29 1.275 0.62 3.075 ;
      RECT 0.095 0.265 0.375 1.82 ;
      RECT 0.095 1.275 1.385 1.535 ;
  END
END scs130lp_clkbuflp_2

MACRO scs130lp_clkbuflp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuflp_4 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.692 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.135 0.715 1.565 ;
        RECT 0.125 1.135 0.41 1.78 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.355 1.17 3.74 1.79 ;
        RECT 2.745 1.17 3.075 3.075 ;
        RECT 2.355 0.325 2.775 1.875 ;
        RECT 1.685 1.705 3.075 1.875 ;
        RECT 2.195 0.325 2.775 0.655 ;
        RECT 1.685 1.705 2.015 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.985 -0.085 3.315 0.655 ;
        RECT 1.405 -0.085 1.735 0.655 ;
        RECT 0.125 -0.085 0.425 0.895 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.275 2.085 3.605 3.415 ;
        RECT 2.215 2.085 2.545 3.415 ;
        RECT 1.225 2.065 1.485 3.415 ;
        RECT 0.125 2.065 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.625 2.065 1.055 3.075 ;
      RECT 0.885 0.255 1.055 3.075 ;
      RECT 0.885 1.205 2.13 1.535 ;
      RECT 0.885 0.255 1.23 1.535 ;
  END
END scs130lp_clkbuflp_4

MACRO scs130lp_clkbuflp_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkbuflp_8 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.384 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.14 0.715 1.565 ;
        RECT 0.125 1.14 0.425 1.88 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.428 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.875 0.265 6.735 1.79 ;
        RECT 5.925 0.265 6.255 3.075 ;
        RECT 4.1 1.17 6.735 1.79 ;
        RECT 4.865 1.17 5.195 3.075 ;
        RECT 4.1 0.775 4.96 1.875 ;
        RECT 4.585 0.345 4.96 1.875 ;
        RECT 3.805 1.705 4.135 3.075 ;
        RECT 3.005 0.775 4.96 1.035 ;
        RECT 2.745 1.705 4.135 1.885 ;
        RECT 3.005 0.345 3.335 1.035 ;
        RECT 2.745 1.705 3.075 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 5.375 -0.085 5.705 0.675 ;
        RECT 3.795 -0.085 4.125 0.605 ;
        RECT 1.675 -0.085 2.55 0.875 ;
        RECT 0.125 -0.085 0.425 0.89 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.455 2.085 6.785 3.415 ;
        RECT 5.395 2.085 5.725 3.415 ;
        RECT 4.335 2.085 4.665 3.415 ;
        RECT 3.275 2.085 3.605 3.415 ;
        RECT 2.215 2.085 2.545 3.415 ;
        RECT 1.155 2.11 1.485 3.415 ;
        RECT 0.095 2.065 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.66 1.205 1.995 3.075 ;
      RECT 0.625 1.77 0.955 3.075 ;
      RECT 0.955 1.205 1.995 1.94 ;
      RECT 0.955 1.205 3.87 1.535 ;
      RECT 0.955 0.255 1.23 1.94 ;
      RECT 0.885 0.255 1.23 0.985 ;
  END
END scs130lp_clkbuflp_8

MACRO scs130lp_clkdlybuf4s15_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s15_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s15_1

MACRO scs130lp_clkdlybuf4s15_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s15_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.875 1.815 4.125 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s15_2

MACRO scs130lp_clkdlybuf4s18_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s18_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s18_1

MACRO scs130lp_clkdlybuf4s18_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s18_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.875 1.815 4.125 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s18_2

MACRO scs130lp_clkdlybuf4s25_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s25_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s25_1

MACRO scs130lp_clkdlybuf4s25_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s25_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.875 1.815 4.125 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s25_2

MACRO scs130lp_clkdlybuf4s50_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s50_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s50_1

MACRO scs130lp_clkdlybuf4s50_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkdlybuf4s50_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.875 1.815 4.125 3.415 ;
        RECT 2.71 2.165 3.04 3.415 ;
        RECT 0.595 2.38 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_clkdlybuf4s50_2

MACRO scs130lp_clkinv_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_0 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.4 2.13 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 0.78 0.875 2.96 ;
        RECT 0.605 0.395 0.875 2.96 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
        RECT 0.105 -0.085 0.435 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
        RECT 0.105 2.3 0.4 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_0

MACRO scs130lp_clkinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.79 0.475 1.8 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.645 0.84 1.285 1.9 ;
        RECT 0.645 0.84 0.875 2.97 ;
        RECT 0.645 0.395 0.845 2.97 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 1.015 -0.085 1.345 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 1.045 2.18 1.345 3.415 ;
        RECT 0.155 2.18 0.475 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_1

MACRO scs130lp_clkinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_16 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 5.544 LAYER li ;
      ANTENNAGATEAREA 5.544 LAYER met1 ;
      ANTENNAMAXAREACAR 0.136296 LAYER li ;
      ANTENNAMAXAREACAR 0.136296 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.075397 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.075397 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.020851 LAYER mcon ;
    PORT
      LAYER li ;
        RECT 8.92 1.16 10.545 1.625 ;
        RECT 8.06 1.16 8.325 1.625 ;
        RECT 7.2 1.16 7.465 1.625 ;
        RECT 6.34 1.16 6.605 1.625 ;
        RECT 5.48 1.16 5.745 1.625 ;
        RECT 4.62 1.16 4.885 1.625 ;
        RECT 3.76 1.16 4.025 1.625 ;
        RECT 2.9 1.16 3.165 1.625 ;
        RECT 0.59 1.16 2.305 1.625 ;
      LAYER met1 ;
        RECT 0.715 1.18 10.525 1.41 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3528 LAYER li ;
    ANTENNADIFFAREA 5.1744 LAYER met1 ;
    PORT
      LAYER li ;
        RECT 10.21 1.835 10.47 3.055 ;
        RECT 9.355 1.835 9.61 3.055 ;
        RECT 8.495 0.395 8.75 3.055 ;
        RECT 7.635 0.395 7.89 3.055 ;
        RECT 6.775 0.395 7.03 3.055 ;
        RECT 5.915 0.395 6.17 3.055 ;
        RECT 5.05 1.885 5.31 3.055 ;
        RECT 5.055 0.395 5.31 3.055 ;
        RECT 4.195 0.395 4.45 3.055 ;
        RECT 3.335 0.395 3.59 3.055 ;
        RECT 2.475 0.395 2.73 3.055 ;
        RECT 1.615 1.835 1.87 3.055 ;
        RECT 0.755 1.835 1.01 3.055 ;
      LAYER met1 ;
        RECT 0.735 1.92 10.485 2.15 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 8.92 -0.085 9.185 0.725 ;
        RECT 8.06 -0.085 8.325 0.725 ;
        RECT 7.2 -0.085 7.465 0.725 ;
        RECT 6.34 -0.085 6.605 0.725 ;
        RECT 5.48 -0.085 5.745 0.725 ;
        RECT 4.62 -0.085 4.885 0.725 ;
        RECT 3.76 -0.085 4.025 0.725 ;
        RECT 2.9 -0.085 3.165 0.725 ;
        RECT 2.035 -0.085 2.305 0.725 ;
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 11.04 3.415 ;
        RECT 10.64 1.835 10.895 3.415 ;
        RECT 9.78 1.835 10.04 3.415 ;
        RECT 8.92 1.835 9.18 3.415 ;
        RECT 8.06 1.835 8.32 3.415 ;
        RECT 7.2 1.835 7.46 3.415 ;
        RECT 6.34 1.835 6.6 3.415 ;
        RECT 5.48 1.835 5.74 3.415 ;
        RECT 4.62 1.835 4.88 3.415 ;
        RECT 3.76 1.835 4.02 3.415 ;
        RECT 2.9 1.835 3.16 3.415 ;
        RECT 2.04 1.835 2.3 3.415 ;
        RECT 1.18 1.835 1.44 3.415 ;
        RECT 0.32 1.835 0.58 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_16

MACRO scs130lp_clkinv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_2 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.693 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.415 1.21 1.425 1.545 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8043 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.715 1.78 1.885 ;
        RECT 1.595 0.84 1.78 1.885 ;
        RECT 1.1 0.84 1.78 1.04 ;
        RECT 1.1 0.395 1.325 1.04 ;
        RECT 1.01 1.715 1.27 3.045 ;
        RECT 0.155 1.715 0.41 3.045 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.495 -0.085 1.825 0.67 ;
        RECT 0.635 -0.085 0.93 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.44 2.055 1.695 3.415 ;
        RECT 0.58 2.055 0.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_2

MACRO scs130lp_clkinv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_4 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.386 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 1.21 2.865 1.545 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.23 1.715 3.22 1.885 ;
        RECT 3.035 0.84 3.22 1.885 ;
        RECT 0.23 0.84 3.22 1.04 ;
        RECT 2.45 1.715 2.71 3.045 ;
        RECT 2.02 0.395 2.275 1.04 ;
        RECT 1.595 1.715 1.85 3.045 ;
        RECT 1.16 0.395 1.42 1.04 ;
        RECT 0.735 1.715 0.99 3.045 ;
        RECT 0.23 0.84 0.4 1.885 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.445 -0.085 2.745 0.67 ;
        RECT 1.59 -0.085 1.85 0.67 ;
        RECT 0.695 -0.085 0.99 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.88 2.055 3.135 3.415 ;
        RECT 2.02 2.055 2.28 3.415 ;
        RECT 1.16 2.055 1.42 3.415 ;
        RECT 0.3 2.055 0.56 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_4

MACRO scs130lp_clkinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_8 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.772 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.515 1.21 5.265 1.54 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.175 1.71 5.62 1.885 ;
        RECT 5.435 0.84 5.62 1.885 ;
        RECT 0.175 0.84 5.62 1.04 ;
        RECT 4.93 1.71 5.19 3.045 ;
        RECT 4.075 1.71 4.33 3.045 ;
        RECT 4.07 0.395 4.33 1.04 ;
        RECT 3.215 1.71 3.47 3.045 ;
        RECT 3.21 0.395 3.47 1.04 ;
        RECT 2.355 1.71 2.61 3.045 ;
        RECT 2.35 0.395 2.61 1.04 ;
        RECT 1.495 1.71 1.75 3.045 ;
        RECT 1.49 0.395 1.75 1.04 ;
        RECT 0.635 1.71 0.89 3.045 ;
        RECT 0.175 0.84 0.345 1.885 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.5 -0.085 4.795 0.67 ;
        RECT 3.64 -0.085 3.9 0.67 ;
        RECT 2.78 -0.085 3.04 0.67 ;
        RECT 1.92 -0.085 2.18 0.67 ;
        RECT 1.025 -0.085 1.32 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.36 2.055 5.615 3.415 ;
        RECT 4.5 2.055 4.76 3.415 ;
        RECT 3.64 2.055 3.9 3.415 ;
        RECT 2.78 2.055 3.04 3.415 ;
        RECT 1.92 2.055 2.18 3.415 ;
        RECT 1.06 2.055 1.32 3.415 ;
        RECT 0.2 2.055 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_8

MACRO scs130lp_clkinv_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_lp 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 2.15 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3021 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 2.32 1.315 3 ;
        RECT 1.085 0.44 1.315 3 ;
        RECT 0.985 0.44 1.315 0.9 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.165 -0.085 0.495 0.9 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.165 2.32 0.495 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_lp

MACRO scs130lp_clkinv_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinv_lp2 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.955 0.835 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.96 1.315 3 ;
        RECT 1.085 0.315 1.315 3 ;
        RECT 0.985 0.315 1.315 0.775 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.165 -0.085 0.495 0.775 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.455 1.96 0.785 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinv_lp2

MACRO scs130lp_clkinvlp_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinvlp_16 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 5.65 LAYER li ;
      ANTENNAGATEAREA 5.65 LAYER met1 ;
      ANTENNAMAXAREACAR 0.068823 LAYER li ;
      ANTENNAMAXAREACAR 0.068823 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.049381 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.049381 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.01023 LAYER mcon ;
    PORT
      LAYER li ;
        RECT 7.705 1.18 8.715 1.565 ;
        RECT 6.37 1.18 6.7 1.565 ;
        RECT 4.655 1.18 5.38 1.565 ;
        RECT 3.275 1.18 3.71 1.565 ;
        RECT 1.075 1.18 2.265 1.565 ;
        RECT 0.1 1.105 0.455 1.78 ;
      LAYER met1 ;
        RECT 0.075 1.18 8.545 1.41 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.28 LAYER li ;
    ANTENNADIFFAREA 3.01 LAYER met1 ;
    PORT
      LAYER li ;
        RECT 8.045 1.92 8.375 3 ;
        RECT 7.205 0.445 7.535 1.565 ;
        RECT 6.985 1.195 7.315 3 ;
        RECT 5.895 1.875 6.255 3 ;
        RECT 5.895 1.195 6.19 3 ;
        RECT 5.625 0.445 5.955 1.565 ;
        RECT 4.865 1.92 5.195 3 ;
        RECT 4.045 0.445 4.375 1.565 ;
        RECT 3.805 1.805 4.135 3 ;
        RECT 3.88 1.195 4.135 3 ;
        RECT 2.745 1.195 3.075 3 ;
        RECT 2.465 0.445 2.795 1.565 ;
        RECT 1.685 1.92 2.015 3 ;
        RECT 0.625 0.315 1.215 0.78 ;
        RECT 0.625 1.735 0.955 3 ;
        RECT 0.625 0.315 0.955 1.01 ;
        RECT 0.625 0.315 0.905 3 ;
      LAYER met1 ;
        RECT 0.575 1.92 8.355 2.15 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 7.995 -0.085 8.325 0.775 ;
        RECT 6.415 -0.085 6.745 0.775 ;
        RECT 4.835 -0.085 5.165 0.775 ;
        RECT 3.255 -0.085 3.585 0.775 ;
        RECT 1.675 -0.085 2.005 0.775 ;
        RECT 0.095 -0.085 0.425 0.775 ;
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 8.575 1.96 8.905 3.415 ;
        RECT 7.515 1.96 7.845 3.415 ;
        RECT 6.455 1.96 6.785 3.415 ;
        RECT 5.395 1.96 5.725 3.415 ;
        RECT 4.335 1.96 4.665 3.415 ;
        RECT 3.275 1.96 3.605 3.415 ;
        RECT 2.215 1.96 2.545 3.415 ;
        RECT 1.155 1.96 1.485 3.415 ;
        RECT 0.095 1.96 0.425 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinvlp_16

MACRO scs130lp_clkinvlp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinvlp_2 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.665 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 0.995 0.855 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 0.315 1.62 0.78 ;
        RECT 0.93 1.96 1.32 3 ;
        RECT 1.035 0.315 1.32 3 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.47 -0.085 0.8 0.775 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.49 1.96 1.79 3.415 ;
        RECT 0.4 1.96 0.73 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinvlp_2

MACRO scs130lp_clkinvlp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinvlp_4 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.33 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.105 0.455 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.685 1.235 2.015 3 ;
        RECT 0.625 1.235 2.015 1.565 ;
        RECT 0.625 0.315 1.215 0.78 ;
        RECT 0.625 0.315 0.955 3 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.675 -0.085 2.005 0.775 ;
        RECT 0.095 -0.085 0.425 0.775 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.215 1.96 2.545 3.415 ;
        RECT 1.155 1.96 1.485 3.415 ;
        RECT 0.095 1.96 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinvlp_4

MACRO scs130lp_clkinvlp_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_clkinvlp_8 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.66 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.105 0.455 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.428 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.805 1.195 4.135 3 ;
        RECT 0.625 1.195 4.135 1.565 ;
        RECT 2.745 1.195 3.075 3 ;
        RECT 2.465 0.445 2.795 1.565 ;
        RECT 1.685 1.195 2.015 3 ;
        RECT 0.625 0.315 1.215 0.78 ;
        RECT 0.625 0.315 0.955 3 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.255 -0.085 3.585 0.775 ;
        RECT 1.675 -0.085 2.005 0.775 ;
        RECT 0.095 -0.085 0.425 0.775 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.335 1.96 4.665 3.415 ;
        RECT 3.275 1.96 3.605 3.415 ;
        RECT 2.215 1.96 2.545 3.415 ;
        RECT 1.155 1.96 1.485 3.415 ;
        RECT 0.095 1.96 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_clkinvlp_8

MACRO scs130lp_conb_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_conb_0 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1792 LAYER li ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.18 0.865 2.97 ;
        RECT 0.28 1.18 0.865 2.12 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1176 LAYER li ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 0.84 1.355 2.12 ;
        RECT 0.62 0.84 1.355 1.01 ;
        RECT 0.62 0.46 0.845 1.01 ;
    END
  END LO
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 1.015 -0.085 1.345 0.67 ;
        RECT 0.155 -0.085 0.45 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 1.035 2.29 1.345 3.415 ;
        RECT 0.155 2.29 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_conb_0

MACRO scs130lp_conb_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_conb_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1792 LAYER li ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.18 0.855 2.97 ;
        RECT 0.28 1.18 0.855 2.12 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1176 LAYER li ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 0.84 1.355 2.12 ;
        RECT 0.62 0.84 1.355 1.01 ;
        RECT 0.62 0.395 0.845 1.01 ;
    END
  END LO
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 1.015 -0.085 1.345 0.67 ;
        RECT 0.155 -0.085 0.45 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 1.025 2.29 1.345 3.415 ;
        RECT 0.155 2.29 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_conb_1

MACRO scs130lp_decap_12
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decap_12 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.93 -0.085 5.26 1.125 ;
        RECT 0.65 1.605 2.58 1.935 ;
        RECT 0.65 -0.085 0.98 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.865 1.34 5.195 3.415 ;
        RECT 2.925 1.34 5.195 1.675 ;
        RECT 0.575 2.105 0.905 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decap_12

MACRO scs130lp_decap_3
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decap_3 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.95 -0.085 1.28 0.625 ;
        RECT 0.17 1.605 0.66 1.935 ;
        RECT 0.17 -0.085 0.5 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.885 0.86 1.215 3.415 ;
        RECT 0.67 0.86 1.215 1.225 ;
        RECT 0.095 2.105 0.425 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decap_3

MACRO scs130lp_decap_4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decap_4 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.45 -0.085 1.78 1.125 ;
        RECT 0.17 1.605 0.74 1.935 ;
        RECT 0.17 -0.085 0.5 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.385 1.34 1.715 3.415 ;
        RECT 1.18 1.34 1.715 1.675 ;
        RECT 0.095 2.105 0.425 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decap_4

MACRO scs130lp_decap_6
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decap_6 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.45 -0.085 2.78 1.17 ;
        RECT 0.17 1.605 1.08 1.935 ;
        RECT 0.17 -0.085 0.5 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.385 1.34 2.715 3.415 ;
        RECT 1.555 1.34 2.715 1.675 ;
        RECT 0.095 2.105 0.425 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decap_6

MACRO scs130lp_decap_8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decap_8 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.93 -0.085 3.26 1.125 ;
        RECT 0.65 1.605 1.56 1.935 ;
        RECT 0.65 -0.085 0.98 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.865 1.34 3.195 3.415 ;
        RECT 1.955 1.34 3.195 1.675 ;
        RECT 0.575 2.105 0.905 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decap_8

MACRO scs130lp_decapkapwr_12
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decapkapwr_12 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 4.865 1.34 5.195 3.075 ;
        RECT 0.575 2.675 5.195 2.945 ;
        RECT 2.925 1.34 5.195 1.675 ;
        RECT 0.575 2.105 0.905 3.075 ;
      LAYER met1 ;
        RECT 0.07 2.675 5.69 2.945 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.93 -0.085 5.26 1.125 ;
        RECT 0.65 1.605 2.58 1.935 ;
        RECT 0.65 -0.085 0.98 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decapkapwr_12

MACRO scs130lp_decapkapwr_3
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decapkapwr_3 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.885 0.86 1.215 3.075 ;
        RECT 0.095 2.675 1.215 2.945 ;
        RECT 0.67 0.86 1.215 1.225 ;
        RECT 0.095 2.105 0.425 3.075 ;
      LAYER met1 ;
        RECT 0.07 2.675 1.37 2.945 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.95 -0.085 1.28 0.625 ;
        RECT 0.17 1.605 0.66 1.935 ;
        RECT 0.17 -0.085 0.5 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decapkapwr_3

MACRO scs130lp_decapkapwr_4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decapkapwr_4 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 1.385 1.34 1.79 3.075 ;
        RECT 0.095 2.675 1.79 2.945 ;
        RECT 1.18 1.34 1.79 1.675 ;
        RECT 0.095 2.105 0.425 3.075 ;
      LAYER met1 ;
        RECT 0.07 2.675 1.85 2.945 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.45 -0.085 1.78 1.125 ;
        RECT 0.17 1.605 0.74 1.935 ;
        RECT 0.17 -0.085 0.5 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decapkapwr_4

MACRO scs130lp_decapkapwr_6
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decapkapwr_6 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 2.385 1.34 2.75 3.075 ;
        RECT 0.095 2.675 2.75 2.945 ;
        RECT 1.555 1.34 2.75 1.675 ;
        RECT 0.095 2.105 0.425 3.075 ;
      LAYER met1 ;
        RECT 0.07 2.675 2.81 2.945 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.45 -0.085 2.78 1.17 ;
        RECT 0.17 1.605 1.08 1.935 ;
        RECT 0.17 -0.085 0.5 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decapkapwr_6

MACRO scs130lp_decapkapwr_8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_decapkapwr_8 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 2.865 1.34 3.285 3.075 ;
        RECT 0.495 2.675 3.285 2.945 ;
        RECT 1.955 1.34 3.285 1.675 ;
        RECT 0.495 2.105 0.905 3.075 ;
      LAYER met1 ;
        RECT 0.07 2.675 3.77 2.945 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.93 -0.085 3.26 1.125 ;
        RECT 0.65 1.605 1.56 1.935 ;
        RECT 0.65 -0.085 0.98 1.935 ;
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_decapkapwr_8

MACRO scs130lp_dfbbn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfbbn_1 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 0.955 0.445 2.15 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.18 2.08 1.51 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.475 1.815 13.83 3.065 ;
        RECT 13.66 0.265 13.83 3.065 ;
        RECT 13.475 0.265 13.83 1.125 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5859 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.075 1.695 12.435 2.995 ;
        RECT 12.265 0.265 12.435 2.995 ;
        RECT 11.975 0.265 12.435 1.005 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.165 1.18 11.52 1.515 ;
    END
  END RESETB
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 1.166892 LAYER li ;
      ANTENNAMAXAREACAR 1.166892 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.004505 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.004505 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 8.735 1.55 9.025 1.78 ;
        RECT 4.895 1.595 9.025 1.735 ;
        RECT 4.895 1.55 5.185 1.78 ;
      LAYER li ;
        RECT 8.795 1.5 9.58 1.83 ;
        RECT 4.875 1.405 5.155 1.78 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.92 0.085 ;
        RECT 13.045 -0.085 13.295 1.125 ;
        RECT 11.545 -0.085 11.795 1 ;
        RECT 8.945 -0.085 9.275 0.97 ;
        RECT 6.835 -0.085 7.085 0.905 ;
        RECT 4.18 -0.085 4.51 0.875 ;
        RECT 1.595 -0.085 1.925 1 ;
        RECT 0.11 -0.085 0.36 0.775 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.92 3.415 ;
        RECT 13.045 1.815 13.295 3.415 ;
        RECT 11.565 2.555 11.895 3.415 ;
        RECT 10.515 2.555 10.845 3.415 ;
        RECT 9.215 2.58 9.545 3.415 ;
        RECT 6.725 1.875 7.055 3.415 ;
        RECT 4.605 2.66 4.935 3.415 ;
        RECT 1.715 2.225 2.045 3.415 ;
        RECT 0.115 2.385 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 12.615 0.665 12.865 2.495 ;
      RECT 12.615 1.305 13.48 1.635 ;
      RECT 9.725 2.07 10.055 3.065 ;
      RECT 8.86 2.07 10.055 2.4 ;
      RECT 8.86 2.205 11.895 2.375 ;
      RECT 11.725 1.185 11.895 2.375 ;
      RECT 10.3 0.83 10.47 2.375 ;
      RECT 11.725 1.185 12.085 1.515 ;
      RECT 10.125 0.83 10.47 1 ;
      RECT 9.965 0.615 10.295 0.97 ;
      RECT 10.65 1.695 11.39 2.025 ;
      RECT 10.65 0.83 10.98 2.025 ;
      RECT 10.65 0.83 11.365 1 ;
      RECT 11.035 0.635 11.365 1 ;
      RECT 9.455 0.265 9.785 0.97 ;
      RECT 10.475 0.265 10.805 0.65 ;
      RECT 9.455 0.265 10.805 0.435 ;
      RECT 7.71 2.12 8.1 2.715 ;
      RECT 7.93 0.575 8.1 2.715 ;
      RECT 9.775 1.46 10.12 1.79 ;
      RECT 9.775 1.15 9.945 1.79 ;
      RECT 7.93 1.15 9.945 1.32 ;
      RECT 7.93 0.575 8.26 1.32 ;
      RECT 7.36 2.895 8.615 3.065 ;
      RECT 8.32 1.73 8.615 3.065 ;
      RECT 7.36 1.085 7.53 3.065 ;
      RECT 3.43 1.055 3.62 1.75 ;
      RECT 7.36 1.345 7.75 1.675 ;
      RECT 6.485 1.085 7.53 1.255 ;
      RECT 3.43 1.055 4.86 1.225 ;
      RECT 4.69 0.265 4.86 1.225 ;
      RECT 6.485 0.265 6.655 1.255 ;
      RECT 4.69 0.265 6.655 0.435 ;
      RECT 5.685 1.915 6.015 2.755 ;
      RECT 4.15 2.31 6.015 2.48 ;
      RECT 4.15 1.755 4.345 2.48 ;
      RECT 5.685 1.915 6.545 2.085 ;
      RECT 6.375 1.435 6.545 2.085 ;
      RECT 6.135 1.435 7.18 1.695 ;
      RECT 6.135 1.125 6.305 1.695 ;
      RECT 5.55 1.125 6.305 1.295 ;
      RECT 5.55 0.965 5.88 1.295 ;
      RECT 5.04 0.615 5.37 0.99 ;
      RECT 6.135 0.615 6.305 0.945 ;
      RECT 5.04 0.615 6.305 0.785 ;
      RECT 3.08 2.225 3.41 2.685 ;
      RECT 3.08 2.225 3.97 2.395 ;
      RECT 3.8 1.405 3.97 2.395 ;
      RECT 3.08 0.53 3.25 2.685 ;
      RECT 4.525 1.96 5.505 2.13 ;
      RECT 5.335 1.475 5.505 2.13 ;
      RECT 4.525 1.405 4.695 2.13 ;
      RECT 5.335 1.475 5.955 1.735 ;
      RECT 3.8 1.405 4.695 1.575 ;
      RECT 2.92 0.53 3.25 0.95 ;
      RECT 2.275 2.305 2.605 2.685 ;
      RECT 2.275 2.305 2.9 2.475 ;
      RECT 2.73 1.13 2.9 2.475 ;
      RECT 2.41 0.575 2.74 1.3 ;
      RECT 1.205 2.045 1.535 2.905 ;
      RECT 2.29 1.48 2.55 2.045 ;
      RECT 1.245 1.875 2.55 2.045 ;
      RECT 1.245 0.575 1.415 2.905 ;
      RECT 1.085 0.575 1.415 1.015 ;
      RECT 0.625 1.195 0.955 3.065 ;
      RECT 0.625 1.195 1.065 1.865 ;
      RECT 0.625 0.315 0.87 3.065 ;
      RECT 0.54 0.315 0.87 0.775 ;
  END
END scs130lp_dfbbn_1

MACRO scs130lp_dfbbn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfbbn_2 0 0 ;
  SIZE 14.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.91 0.435 2.15 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.18 2.085 1.51 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.275 0.925 14.445 1.955 ;
        RECT 14.01 1.785 14.34 3.065 ;
        RECT 14.01 0.265 14.34 1.095 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.15 1.695 12.41 2.99 ;
        RECT 12.24 0.265 12.41 2.99 ;
        RECT 12.08 0.265 12.41 1.005 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.165 1.18 11.56 1.51 ;
    END
  END RESETB
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 1.159459 LAYER li ;
      ANTENNAMAXAREACAR 1.159459 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 8.735 1.55 9.025 1.78 ;
        RECT 4.895 1.595 9.025 1.735 ;
        RECT 4.895 1.55 5.185 1.78 ;
      LAYER li ;
        RECT 8.795 1.47 9.575 1.8 ;
        RECT 4.9 1.405 5.165 1.78 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 14.88 0.085 ;
        RECT 14.52 -0.085 14.77 0.745 ;
        RECT 13.58 -0.085 13.83 1.095 ;
        RECT 12.59 -0.085 12.84 1.095 ;
        RECT 11.65 -0.085 11.9 1 ;
        RECT 9.035 -0.085 9.365 0.94 ;
        RECT 6.86 -0.085 7.11 0.905 ;
        RECT 4.205 -0.085 4.535 0.875 ;
        RECT 1.6 -0.085 1.93 1 ;
        RECT 0.11 -0.085 0.36 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 14.88 3.415 ;
        RECT 14.52 2.135 14.77 3.415 ;
        RECT 13.58 1.815 13.83 3.415 ;
        RECT 12.59 1.69 12.84 3.415 ;
        RECT 11.64 2.55 11.97 3.415 ;
        RECT 10.575 2.55 10.905 3.415 ;
        RECT 9.355 2.55 9.605 3.415 ;
        RECT 6.235 1.875 6.565 3.415 ;
        RECT 4.63 2.66 4.96 3.415 ;
        RECT 1.72 2.225 2.05 3.415 ;
        RECT 0.14 2.385 0.47 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 13.07 0.635 13.4 2.495 ;
      RECT 13.07 1.275 14.095 1.605 ;
      RECT 9.785 2.2 10.115 3 ;
      RECT 8.885 2.2 11.965 2.37 ;
      RECT 11.795 1.185 11.965 2.37 ;
      RECT 10.305 0.615 10.475 2.37 ;
      RECT 8.885 2.04 9.215 2.37 ;
      RECT 11.795 1.185 12.06 1.515 ;
      RECT 10.135 0.615 10.475 1.165 ;
      RECT 10.815 1.69 11.46 2.02 ;
      RECT 10.655 0.83 10.985 1.69 ;
      RECT 10.655 0.83 11.47 1 ;
      RECT 11.22 0.265 11.47 1 ;
      RECT 9.545 0.265 9.875 0.94 ;
      RECT 10.655 0.265 10.905 0.65 ;
      RECT 9.545 0.265 10.905 0.435 ;
      RECT 7.685 2.12 8.125 2.715 ;
      RECT 7.955 0.575 8.125 2.715 ;
      RECT 9.785 1.345 10.125 1.675 ;
      RECT 9.785 1.12 9.955 1.675 ;
      RECT 7.955 1.12 9.955 1.29 ;
      RECT 7.955 0.575 8.285 1.29 ;
      RECT 7.335 2.895 8.615 3.065 ;
      RECT 8.345 1.7 8.615 3.065 ;
      RECT 7.335 1.085 7.505 3.065 ;
      RECT 3.44 1.055 3.64 1.76 ;
      RECT 7.335 1.085 7.775 1.675 ;
      RECT 6.51 1.085 7.775 1.255 ;
      RECT 3.44 1.055 4.885 1.225 ;
      RECT 4.715 0.265 4.885 1.225 ;
      RECT 6.51 0.265 6.68 1.255 ;
      RECT 4.715 0.265 6.68 0.435 ;
      RECT 5.14 2.31 5.47 2.755 ;
      RECT 4.17 2.31 6.055 2.48 ;
      RECT 5.885 1.125 6.055 2.48 ;
      RECT 4.17 1.755 4.37 2.48 ;
      RECT 6.825 1.435 7.155 1.735 ;
      RECT 5.885 1.435 7.155 1.605 ;
      RECT 5.575 0.965 5.905 1.295 ;
      RECT 5.065 0.615 5.395 0.96 ;
      RECT 6.16 0.615 6.33 0.945 ;
      RECT 5.065 0.615 6.33 0.785 ;
      RECT 3.09 2.225 3.42 2.685 ;
      RECT 3.09 2.225 3.99 2.395 ;
      RECT 3.82 1.405 3.99 2.395 ;
      RECT 3.09 0.5 3.26 2.685 ;
      RECT 4.55 1.96 5.705 2.13 ;
      RECT 5.375 1.475 5.705 2.13 ;
      RECT 4.55 1.405 4.72 2.13 ;
      RECT 3.82 1.405 4.72 1.575 ;
      RECT 3.035 0.5 3.26 0.95 ;
      RECT 2.29 2.305 2.62 2.685 ;
      RECT 2.29 2.305 2.91 2.475 ;
      RECT 2.74 1.13 2.91 2.475 ;
      RECT 2.445 0.575 2.775 1.3 ;
      RECT 1.21 1.875 1.54 2.905 ;
      RECT 1.21 1.875 2.56 2.045 ;
      RECT 2.295 1.48 2.56 2.045 ;
      RECT 1.21 0.575 1.38 2.905 ;
      RECT 1.09 0.575 1.42 1 ;
      RECT 0.65 1.3 1.005 3.065 ;
      RECT 0.65 0.265 0.87 3.065 ;
      RECT 0.54 0.265 0.87 0.725 ;
  END
END scs130lp_dfbbn_2

MACRO scs130lp_dfbbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfbbp_1 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.905 0.455 2.15 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.77 0.765 2.28 2.055 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.505 1.815 12.87 3.065 ;
        RECT 12.7 0.265 12.87 3.065 ;
        RECT 12.505 0.265 12.87 1.095 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.085 1.695 11.445 2.995 ;
        RECT 11.275 0.265 11.445 2.995 ;
        RECT 11.01 0.265 11.445 1.005 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.205 1.18 10.55 1.515 ;
    END
  END RESETB
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 1.057432 LAYER li ;
      ANTENNAMAXAREACAR 1.057432 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.968468 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.968468 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 8.255 1.92 8.545 2.15 ;
        RECT 4.415 1.965 8.545 2.105 ;
        RECT 4.415 1.92 4.705 2.15 ;
      LAYER li ;
        RECT 8.265 1.66 8.56 2.15 ;
        RECT 4.375 1.405 4.705 1.78 ;
        RECT 4.375 1.405 4.675 2.15 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.96 0.085 ;
        RECT 12.075 -0.085 12.325 0.935 ;
        RECT 10.58 -0.085 10.83 1 ;
        RECT 8.07 -0.085 8.32 0.765 ;
        RECT 6.14 -0.085 6.39 0.58 ;
        RECT 4.05 -0.085 4.38 0.875 ;
        RECT 1.765 -0.085 2.095 0.585 ;
        RECT 0.115 -0.085 0.365 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.96 3.415 ;
        RECT 12.075 1.815 12.325 3.415 ;
        RECT 10.575 2.555 10.905 3.415 ;
        RECT 9.5 2.555 9.83 3.415 ;
        RECT 8.14 2.68 8.47 3.415 ;
        RECT 5.595 2.31 5.925 3.415 ;
        RECT 4.265 2.68 4.595 3.415 ;
        RECT 1.765 2.585 2.095 3.415 ;
        RECT 0.185 2.385 0.515 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 6.815 1.18 7.105 1.41 ;
      RECT 2.495 1.18 2.785 1.41 ;
      RECT 2.495 1.225 7.105 1.365 ;
    LAYER li ;
      RECT 11.645 1.465 11.895 2.495 ;
      RECT 11.645 1.465 12.52 1.635 ;
      RECT 12.155 1.305 12.52 1.635 ;
      RECT 12.155 1.115 12.325 1.635 ;
      RECT 11.645 1.115 12.325 1.285 ;
      RECT 11.645 0.635 11.895 1.285 ;
      RECT 8.74 2.145 8.99 3.01 ;
      RECT 7.765 2.33 8.99 2.5 ;
      RECT 10.735 1.185 10.905 2.375 ;
      RECT 8.74 2.205 10.905 2.375 ;
      RECT 7.765 1.66 8.055 2.5 ;
      RECT 8.74 2.145 9.485 2.375 ;
      RECT 9.315 1.125 9.485 2.375 ;
      RECT 10.735 1.185 11.095 1.515 ;
      RECT 9.09 1.125 9.485 1.455 ;
      RECT 9.68 1.695 10.395 2.025 ;
      RECT 9.68 0.775 10.01 2.025 ;
      RECT 5.73 0.76 6.015 1.315 ;
      RECT 7.665 0.945 8.91 1.115 ;
      RECT 9.68 0.775 10.4 1 ;
      RECT 10.07 0.635 10.4 1 ;
      RECT 8.74 0.775 10.4 0.945 ;
      RECT 7.665 0.265 7.835 1.115 ;
      RECT 5.73 0.76 6.74 0.93 ;
      RECT 6.57 0.265 6.74 0.93 ;
      RECT 6.57 0.265 7.835 0.435 ;
      RECT 6.64 2.58 6.97 3 ;
      RECT 6.64 2.58 7.585 2.75 ;
      RECT 7.415 1.31 7.585 2.75 ;
      RECT 8.74 1.635 9.135 1.965 ;
      RECT 8.74 1.31 8.91 1.965 ;
      RECT 7.315 1.31 8.91 1.48 ;
      RECT 7.315 0.615 7.485 1.48 ;
      RECT 6.96 0.615 7.485 0.93 ;
      RECT 6.805 2.07 7.235 2.4 ;
      RECT 6.805 1.11 7.135 2.4 ;
      RECT 4.855 1.96 5.105 2.755 ;
      RECT 3.88 2.33 5.105 2.5 ;
      RECT 3.88 1.405 4.165 2.5 ;
      RECT 4.855 1.96 6.555 2.13 ;
      RECT 6.225 1.11 6.555 2.13 ;
      RECT 5.38 0.705 5.55 2.13 ;
      RECT 5.07 0.615 5.4 0.875 ;
      RECT 4.56 0.265 4.89 0.875 ;
      RECT 5.58 0.265 5.91 0.525 ;
      RECT 4.56 0.265 5.91 0.435 ;
      RECT 3.32 2.41 3.7 2.755 ;
      RECT 3.53 0.48 3.7 2.755 ;
      RECT 4.915 1.055 5.2 1.385 ;
      RECT 3.53 1.055 5.2 1.225 ;
      RECT 3.14 0.48 3.7 0.65 ;
      RECT 3.14 0.265 3.47 0.65 ;
      RECT 2.81 2.06 3.14 2.755 ;
      RECT 2.81 2.06 3.35 2.23 ;
      RECT 3.18 0.83 3.35 2.23 ;
      RECT 2.63 0.83 3.35 1 ;
      RECT 2.63 0.265 2.96 1 ;
      RECT 1.255 0.265 1.585 2.975 ;
      RECT 1.255 2.235 2.63 2.405 ;
      RECT 2.46 1.18 2.63 2.405 ;
      RECT 2.46 1.56 3 1.88 ;
      RECT 2.46 1.18 2.755 1.88 ;
      RECT 1.105 0.265 1.585 0.675 ;
      RECT 0.695 1.27 1.025 3.065 ;
      RECT 0.695 0.265 0.875 3.065 ;
      RECT 0.545 0.265 0.875 0.725 ;
      RECT 8.5 0.265 9.845 0.595 ;
  END
END scs130lp_dfbbp_1

MACRO scs130lp_dfrbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfrbp_1 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.53 1.58 0.915 2.18 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 1.39 2.575 2.155 ;
        RECT 2.03 1.21 2.315 2.155 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5733 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.17 1.845 10.43 3.075 ;
        RECT 10.225 0.965 10.43 3.075 ;
        RECT 10.09 0.965 10.43 1.165 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5817 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.035 1.82 11.435 3.075 ;
        RECT 11.185 0.255 11.435 3.075 ;
        RECT 11.165 0.255 11.435 1.095 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.378 LAYER met1 ;
      ANTENNAMAXAREACAR 0.680952 LAYER li ;
      ANTENNAMAXAREACAR 0.680952 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.936508 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.936508 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.92 8.065 2.15 ;
        RECT 1.535 1.965 8.065 2.105 ;
        RECT 4.415 1.92 4.705 2.15 ;
        RECT 1.535 1.92 1.825 2.15 ;
      LAYER li ;
        RECT 7.74 1.94 8.07 2.2 ;
        RECT 4.475 1.79 4.9 2.12 ;
        RECT 1.595 1.45 1.86 2.155 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.52 0.085 ;
        RECT 10.665 -0.085 10.995 0.455 ;
        RECT 9.6 -0.085 9.93 0.455 ;
        RECT 7.495 -0.085 7.685 0.95 ;
        RECT 5.225 -0.085 5.555 0.55 ;
        RECT 1.545 -0.085 1.875 0.7 ;
        RECT 0.6 -0.085 0.81 0.9 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.52 3.415 ;
        RECT 10.6 1.82 10.865 3.415 ;
        RECT 9.505 2.505 9.835 3.415 ;
        RECT 8.59 2.405 8.825 3.415 ;
        RECT 7.325 2.405 7.995 3.415 ;
        RECT 5.35 2.24 5.68 3.415 ;
        RECT 4.34 2.65 4.67 3.415 ;
        RECT 1.97 2.665 2.32 3.415 ;
        RECT 0.53 2.35 0.86 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.5 2.04 6.82 2.915 ;
      RECT 6.62 0.63 6.82 2.915 ;
      RECT 9.345 1.325 9.64 1.995 ;
      RECT 9.46 0.625 9.64 1.995 ;
      RECT 10.825 1.185 11.015 1.515 ;
      RECT 6.62 1.25 8.43 1.43 ;
      RECT 7.875 1.19 8.43 1.43 ;
      RECT 7.875 0.345 8.045 1.43 ;
      RECT 10.825 0.625 10.995 1.515 ;
      RECT 8.96 0.625 10.995 0.795 ;
      RECT 8.96 0.345 9.13 0.795 ;
      RECT 7.875 0.345 9.13 0.515 ;
      RECT 8.995 2.165 9.325 3.065 ;
      RECT 8.995 2.165 10 2.335 ;
      RECT 9.83 1.345 10 2.335 ;
      RECT 8.995 0.965 9.165 3.065 ;
      RECT 9.83 1.345 10.055 1.675 ;
      RECT 8.96 0.965 9.165 1.25 ;
      RECT 8.96 0.965 9.29 1.145 ;
      RECT 8.165 2.345 8.42 2.735 ;
      RECT 8.25 1.6 8.42 2.735 ;
      RECT 7.2 1.6 7.53 2.19 ;
      RECT 8.25 1.6 8.79 1.97 ;
      RECT 8.61 0.685 8.79 1.97 ;
      RECT 7.2 1.6 8.79 1.77 ;
      RECT 8.225 0.685 8.79 1.015 ;
      RECT 1.03 2.35 1.35 3.02 ;
      RECT 1.11 1.58 1.35 3.02 ;
      RECT 1.205 0.87 1.395 2.1 ;
      RECT 3.095 1.615 3.5 1.945 ;
      RECT 6.27 0.72 6.45 1.72 ;
      RECT 3.095 0.63 3.265 1.945 ;
      RECT 1.205 0.87 2.255 1.04 ;
      RECT 2.045 0.63 2.255 1.04 ;
      RECT 0.98 0.585 1.375 0.9 ;
      RECT 4.54 0.72 6.45 0.89 ;
      RECT 2.045 0.63 4.755 0.8 ;
      RECT 5.93 1.9 6.145 2.91 ;
      RECT 5.07 1.9 6.145 2.07 ;
      RECT 4.04 1.44 4.295 2.03 ;
      RECT 5.93 1.06 6.1 2.91 ;
      RECT 5.07 1.44 5.24 2.07 ;
      RECT 4.04 1.44 5.24 1.61 ;
      RECT 5.77 1.06 6.1 1.32 ;
      RECT 4.85 2.3 5.095 2.735 ;
      RECT 3.515 2.37 3.965 2.735 ;
      RECT 3.68 2.3 5.095 2.47 ;
      RECT 3.68 0.97 3.86 2.735 ;
      RECT 5.41 1.06 5.6 1.72 ;
      RECT 3.435 0.97 3.86 1.3 ;
      RECT 3.435 1.06 5.6 1.26 ;
      RECT 3.435 0.97 4.215 1.26 ;
      RECT 2.54 2.325 3.345 2.735 ;
      RECT 2.755 2.3 3.345 2.735 ;
      RECT 1.52 2.325 1.73 2.735 ;
      RECT 1.52 2.325 3.345 2.495 ;
      RECT 2.755 2.115 3.15 2.735 ;
      RECT 2.755 0.98 2.925 2.735 ;
      RECT 2.485 0.98 2.925 1.22 ;
      RECT 0.1 0.585 0.36 3.02 ;
      RECT 0.1 1.07 1.035 1.4 ;
      RECT 0.1 0.585 0.43 1.4 ;
  END
END scs130lp_dfrbp_1

MACRO scs130lp_dfrbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfrbp_2 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 1.495 0.905 2.165 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.06 1.21 2.64 2.155 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.185 0.335 11.41 3.075 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.195 0.82 9.455 2.92 ;
        RECT 9.265 0.255 9.455 2.92 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.378 LAYER met1 ;
      ANTENNAMAXAREACAR 0.759524 LAYER li ;
      ANTENNAMAXAREACAR 0.759524 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.984127 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.984127 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.92 8.065 2.15 ;
        RECT 1.535 1.965 8.065 2.105 ;
        RECT 4.415 1.92 4.705 2.15 ;
        RECT 1.535 1.92 1.825 2.15 ;
      LAYER li ;
        RECT 7.76 1.95 8.05 2.28 ;
        RECT 4.475 1.95 4.92 2.12 ;
        RECT 4.495 1.79 4.92 2.12 ;
        RECT 1.585 1.45 1.89 2.155 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12 0.085 ;
        RECT 11.58 -0.085 11.875 1.205 ;
        RECT 10.66 -0.085 11.015 1.125 ;
        RECT 9.625 -0.085 9.955 1.11 ;
        RECT 8.765 -0.085 9.095 0.65 ;
        RECT 7.455 -0.085 7.785 1.015 ;
        RECT 5.245 -0.085 5.575 0.55 ;
        RECT 1.575 -0.085 1.905 0.7 ;
        RECT 0.57 -0.085 0.83 0.755 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
      LAYER li ;
        RECT 0 3.245 12 3.415 ;
        RECT 11.58 1.815 11.875 3.415 ;
        RECT 10.6 1.815 10.955 3.415 ;
        RECT 9.625 1.62 9.875 3.415 ;
        RECT 8.685 1.94 9.015 3.415 ;
        RECT 7.345 2.525 8.025 3.415 ;
        RECT 5.37 2.24 5.7 3.415 ;
        RECT 4.36 2.65 4.69 3.415 ;
        RECT 1.99 2.665 2.34 3.415 ;
        RECT 0.55 2.335 0.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 10.125 0.385 10.43 2.485 ;
      RECT 10.125 1.295 11.015 1.625 ;
      RECT 10.125 0.385 10.49 1.625 ;
      RECT 8.22 1.6 8.49 2.855 ;
      RECT 7.22 1.6 7.55 2.27 ;
      RECT 7.22 1.6 8.49 1.78 ;
      RECT 7.22 1.6 9.025 1.77 ;
      RECT 8.745 0.82 9.025 1.77 ;
      RECT 8.245 0.82 9.025 1.07 ;
      RECT 6.52 2.04 6.84 2.915 ;
      RECT 6.64 0.63 6.84 2.915 ;
      RECT 6.64 1.24 8.565 1.43 ;
      RECT 1.05 2.335 1.38 3.02 ;
      RECT 1.11 2.305 1.38 3.02 ;
      RECT 1.21 1.935 1.38 3.02 ;
      RECT 1.235 0.87 1.415 2.155 ;
      RECT 3.205 1.615 3.625 1.945 ;
      RECT 6.29 0.72 6.47 1.72 ;
      RECT 3.205 0.63 3.375 1.945 ;
      RECT 1.235 0.87 2.315 1.04 ;
      RECT 2.075 0.63 2.315 1.04 ;
      RECT 4.56 0.72 6.47 0.89 ;
      RECT 1.235 0.395 1.405 2.155 ;
      RECT 2.075 0.63 4.775 0.8 ;
      RECT 1 0.395 1.405 0.755 ;
      RECT 5.95 1.9 6.165 2.91 ;
      RECT 5.09 1.9 6.165 2.07 ;
      RECT 4.135 1.44 4.305 2.03 ;
      RECT 5.95 1.06 6.12 2.91 ;
      RECT 5.09 1.44 5.26 2.07 ;
      RECT 4.135 1.44 5.26 1.61 ;
      RECT 5.79 1.06 6.12 1.32 ;
      RECT 4.87 2.3 5.115 2.735 ;
      RECT 3.535 2.37 3.985 2.735 ;
      RECT 3.795 2.3 5.115 2.47 ;
      RECT 3.795 0.97 3.965 2.735 ;
      RECT 5.43 1.06 5.62 1.72 ;
      RECT 3.545 0.97 3.965 1.3 ;
      RECT 3.545 1.06 5.62 1.26 ;
      RECT 3.545 0.97 4.235 1.26 ;
      RECT 2.56 2.325 3.365 2.735 ;
      RECT 2.81 2.3 3.365 2.735 ;
      RECT 1.55 2.325 1.75 2.735 ;
      RECT 1.55 2.325 3.365 2.495 ;
      RECT 2.81 2.115 3.17 2.735 ;
      RECT 2.81 0.98 3.035 2.735 ;
      RECT 0.12 2.335 0.38 3.02 ;
      RECT 0.12 0.425 0.355 3.02 ;
      RECT 0.12 0.925 1.055 1.255 ;
      RECT 0.12 0.425 0.4 1.255 ;
  END
END scs130lp_dfrbp_2

MACRO scs130lp_dfrbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfrbp_lp 0 0 ;
  SIZE 18.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.565 1.08 14.275 1.41 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.44 2.315 1.46 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 17.785 0.265 18.115 3.065 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.515 0.265 15.845 3.065 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
      ANTENNAGATEAREA 0.567 LAYER met1 ;
      ANTENNAMAXAREACAR 1.169841 LAYER li ;
      ANTENNAMAXAREACAR 1.169841 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.058201 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.058201 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.15291 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 12.095 1.55 12.385 1.78 ;
        RECT 1.055 1.595 12.385 1.735 ;
        RECT 4.895 1.55 5.185 1.78 ;
        RECT 1.055 1.55 1.345 1.78 ;
      LAYER li ;
        RECT 12.125 1.11 12.455 1.78 ;
        RECT 4.925 1.45 5.275 1.78 ;
        RECT 0.985 1.11 1.315 1.78 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 18.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 18.24 0.085 ;
        RECT 16.995 -0.085 17.325 1.125 ;
        RECT 14.49 -0.085 14.82 0.55 ;
        RECT 10.635 -0.085 10.965 0.485 ;
        RECT 6.91 -0.085 7.24 0.995 ;
        RECT 4.715 -0.085 5.045 0.57 ;
        RECT 1.055 -0.085 1.385 0.7 ;
        RECT 1.055 -0.085 1.315 0.94 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 18.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 18.24 3.415 ;
        RECT 16.995 1.815 17.325 3.415 ;
        RECT 14.715 2.29 15.045 3.415 ;
        RECT 12.815 2.66 12.985 3.415 ;
        RECT 10.635 2.655 10.885 3.415 ;
        RECT 6.84 2.395 7.17 3.415 ;
        RECT 4.66 2.66 4.99 3.415 ;
        RECT 1.425 2.66 1.755 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 16.09 0.665 16.42 2.495 ;
      RECT 16.09 1.305 17.605 1.635 ;
      RECT 13.7 1.94 14.03 2.495 ;
      RECT 13.7 1.94 15.335 2.11 ;
      RECT 15.165 0.73 15.335 2.11 ;
      RECT 9.94 0.665 10.27 1.345 ;
      RECT 13.67 0.73 15.335 0.9 ;
      RECT 9.94 0.665 11.315 0.835 ;
      RECT 11.145 0.265 11.315 0.835 ;
      RECT 13.67 0.265 14 0.9 ;
      RECT 11.145 0.265 14 0.435 ;
      RECT 11.415 2.545 12.285 2.715 ;
      RECT 12.115 1.96 12.285 2.715 ;
      RECT 9.075 2.385 10.105 2.715 ;
      RECT 9.935 1.525 10.105 2.715 ;
      RECT 11.415 1.365 11.585 2.715 ;
      RECT 12.115 1.96 13.37 2.13 ;
      RECT 13.04 1.59 13.37 2.13 ;
      RECT 13.04 1.59 14.985 1.76 ;
      RECT 14.725 1.345 14.985 1.76 ;
      RECT 9.43 1.525 11.585 1.695 ;
      RECT 11.215 1.365 11.585 1.695 ;
      RECT 9.43 0.265 9.76 1.695 ;
      RECT 11.065 2.895 12.635 3.065 ;
      RECT 12.465 2.31 12.635 3.065 ;
      RECT 13.165 2.31 13.495 2.99 ;
      RECT 11.065 1.965 11.235 3.065 ;
      RECT 12.465 2.31 13.495 2.48 ;
      RECT 10.905 1.965 11.235 2.425 ;
      RECT 11.765 0.615 11.935 2.365 ;
      RECT 10.51 1.015 10.84 1.345 ;
      RECT 10.51 1.015 11.935 1.185 ;
      RECT 11.765 0.615 13.275 0.865 ;
      RECT 8.62 2.895 10.455 3.065 ;
      RECT 10.285 2.655 10.455 3.065 ;
      RECT 8.62 1.875 8.87 3.065 ;
      RECT 6.05 0.615 6.38 2.725 ;
      RECT 6.05 2.045 8.44 2.215 ;
      RECT 8.27 1.525 8.44 2.215 ;
      RECT 9.08 1.875 9.755 2.205 ;
      RECT 4.375 1.96 6.38 2.13 ;
      RECT 4.375 1.455 4.705 2.13 ;
      RECT 9.08 0.265 9.25 2.205 ;
      RECT 8.27 1.525 9.25 1.695 ;
      RECT 8.92 0.265 9.25 1.695 ;
      RECT 7.815 0.535 8.09 1.865 ;
      RECT 3.515 0.75 3.845 1.46 ;
      RECT 6.56 1.175 8.74 1.345 ;
      RECT 8.41 0.675 8.74 1.345 ;
      RECT 7.815 0.535 8.145 1.345 ;
      RECT 6.56 0.265 6.73 1.345 ;
      RECT 3.515 0.75 5.395 0.92 ;
      RECT 5.225 0.265 5.395 0.92 ;
      RECT 5.225 0.265 6.73 0.435 ;
      RECT 5.52 2.31 5.85 2.725 ;
      RECT 4.025 2.31 5.85 2.48 ;
      RECT 3.165 0.58 3.335 2.365 ;
      RECT 4.025 1.1 4.195 2.48 ;
      RECT 3.165 1.685 4.195 1.855 ;
      RECT 5.54 1.1 5.87 1.77 ;
      RECT 4.025 1.1 5.87 1.27 ;
      RECT 3.005 0.58 3.335 1 ;
      RECT 2.385 2.895 4.385 3.065 ;
      RECT 4.055 2.66 4.385 3.065 ;
      RECT 2.385 2.31 2.635 3.065 ;
      RECT 2.815 2.545 3.845 2.715 ;
      RECT 3.515 2.035 3.845 2.715 ;
      RECT 0.53 1.96 0.86 2.715 ;
      RECT 2.815 1.96 2.985 2.715 ;
      RECT 0.53 1.96 2.985 2.13 ;
      RECT 2.495 0.58 2.825 2.13 ;
      RECT 0.1 2.895 1.21 3.065 ;
      RECT 1.04 2.31 1.21 3.065 ;
      RECT 1.935 2.31 2.185 2.91 ;
      RECT 0.1 2.265 0.35 3.065 ;
      RECT 1.04 2.31 2.185 2.48 ;
  END
END scs130lp_dfrbp_lp

MACRO scs130lp_dfrtn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfrtn_1 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.805 1.57 8.505 2.215 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.15 1.295 1.395 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.145 1.845 10.475 3.075 ;
        RECT 10.205 0.255 10.475 3.075 ;
        RECT 10.155 0.255 10.475 1.09 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.378 LAYER met1 ;
      ANTENNAMAXAREACAR 1.713889 LAYER li ;
      ANTENNAMAXAREACAR 1.713889 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.761905 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.761905 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 6.815 1.55 7.105 1.78 ;
        RECT 0.095 1.595 7.105 1.735 ;
        RECT 2.495 1.55 2.785 1.78 ;
        RECT 0.095 1.55 0.385 1.78 ;
      LAYER li ;
        RECT 7.045 1.58 7.295 2.25 ;
        RECT 6.855 1.58 7.295 1.835 ;
        RECT 2.555 1.565 3.375 1.75 ;
        RECT 0.095 1.565 0.68 2.12 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.725 -0.085 9.985 1.09 ;
        RECT 9.015 0.89 9.215 1.32 ;
        RECT 8.76 0.89 9.215 1.06 ;
        RECT 8.76 -0.085 8.93 1.06 ;
        RECT 6.79 -0.085 7.12 0.71 ;
        RECT 4.47 -0.085 4.8 0.415 ;
        RECT 3.25 -0.085 3.58 0.54 ;
        RECT 0.255 -0.085 0.585 0.98 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.605 1.845 9.975 3.415 ;
        RECT 8.145 2.745 8.335 3.415 ;
        RECT 6.72 2.785 6.92 3.415 ;
        RECT 4.525 2.965 4.855 3.415 ;
        RECT 2.83 2.61 3.16 3.415 ;
        RECT 0.64 2.63 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.12 1.505 9.435 2.495 ;
      RECT 9.385 1.345 10.035 1.675 ;
      RECT 9.385 0.28 9.555 1.675 ;
      RECT 9.18 0.28 9.555 0.61 ;
      RECT 8.505 2.405 8.845 3.075 ;
      RECT 8.675 1.23 8.845 3.075 ;
      RECT 7.09 2.895 7.975 3.065 ;
      RECT 7.805 2.405 7.975 3.065 ;
      RECT 4.025 2.625 4.355 3.065 ;
      RECT 5.2 2.765 6.245 2.935 ;
      RECT 5.92 2.245 6.245 2.935 ;
      RECT 7.09 2.43 7.26 3.065 ;
      RECT 4.025 2.625 5.37 2.795 ;
      RECT 5.92 2.43 7.26 2.6 ;
      RECT 7.805 2.405 8.845 2.575 ;
      RECT 5.92 2.245 6.25 2.6 ;
      RECT 8.215 1.23 8.845 1.4 ;
      RECT 8.215 0.94 8.475 1.4 ;
      RECT 5.54 1.98 5.72 2.585 ;
      RECT 5.54 1.98 5.77 2.155 ;
      RECT 5.54 1.98 5.8 2.115 ;
      RECT 5.54 1.98 5.83 2.1 ;
      RECT 6 0.605 6.17 2.075 ;
      RECT 5.61 1.975 6.17 2.075 ;
      RECT 5.7 1.905 6.17 2.075 ;
      RECT 5.625 1.965 6.17 2.075 ;
      RECT 5.68 1.935 5.72 2.585 ;
      RECT 5.64 1.96 6.17 2.075 ;
      RECT 5.655 1.95 5.72 2.585 ;
      RECT 6 0.88 7.49 1.06 ;
      RECT 7.31 0.265 7.49 1.06 ;
      RECT 6 0.605 6.225 1.06 ;
      RECT 7.31 0.265 8.36 0.49 ;
      RECT 7.465 1.23 7.635 2.725 ;
      RECT 6.515 1.23 6.685 2.05 ;
      RECT 6.515 1.23 7.99 1.4 ;
      RECT 7.66 0.66 7.99 1.4 ;
      RECT 2.155 1.92 4.275 2.1 ;
      RECT 2.155 0.255 2.335 2.1 ;
      RECT 5.385 1.48 5.555 1.81 ;
      RECT 5.385 1.48 5.83 1.735 ;
      RECT 5.66 0.255 5.83 1.735 ;
      RECT 2.155 0.71 4.165 0.88 ;
      RECT 4.97 0.255 5.14 0.765 ;
      RECT 3.915 0.585 5.14 0.765 ;
      RECT 3.915 0.55 4.245 0.765 ;
      RECT 1.47 0.255 2.335 0.48 ;
      RECT 5.66 0.255 6.375 0.435 ;
      RECT 4.97 0.255 6.375 0.425 ;
      RECT 5.025 2.245 5.37 2.455 ;
      RECT 5.025 0.935 5.205 2.455 ;
      RECT 2.505 1.05 2.835 1.395 ;
      RECT 2.505 1.05 4.505 1.22 ;
      RECT 5.025 0.935 5.48 1.205 ;
      RECT 5.31 0.595 5.48 1.205 ;
      RECT 4.335 0.935 5.48 1.105 ;
      RECT 3.33 2.27 3.645 2.735 ;
      RECT 1.735 2.27 2.04 2.735 ;
      RECT 1.735 2.27 4.845 2.44 ;
      RECT 4.675 1.275 4.845 2.44 ;
      RECT 1.735 2.085 1.985 2.735 ;
      RECT 1.805 0.675 1.985 2.735 ;
      RECT 1.16 1.565 1.565 2.735 ;
      RECT 0.1 2.29 0.47 2.735 ;
      RECT 0.1 2.29 1.565 2.46 ;
      RECT 1.465 0.65 1.635 1.82 ;
      RECT 1.15 0.65 1.635 0.98 ;
  END
END scs130lp_dfrtn_1

MACRO scs130lp_dfrtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfrtp_1 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.45 0.47 2.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.97 1.515 2.545 1.84 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.13 1.845 10.475 3.075 ;
        RECT 10.205 0.365 10.475 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.225 1.555 8.145 1.885 ;
        RECT 5.765 2.905 7.395 3.075 ;
        RECT 7.225 1.555 7.395 3.075 ;
        RECT 5.765 2.635 5.935 3.075 ;
        RECT 4.585 2.635 5.935 2.805 ;
        RECT 4.585 2.475 4.915 2.985 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.695 -0.085 10.035 1.165 ;
        RECT 7.51 -0.085 7.84 1.025 ;
        RECT 5.005 -0.085 5.335 0.355 ;
        RECT 2.005 -0.085 2.335 1.005 ;
        RECT 0.595 -0.085 0.785 0.93 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.585 1.845 9.96 3.415 ;
        RECT 8.635 2.63 8.92 3.415 ;
        RECT 7.565 2.63 7.905 3.415 ;
        RECT 5.255 2.975 5.585 3.415 ;
        RECT 3.755 2.795 3.975 3.415 ;
        RECT 1.91 2.845 2.24 3.415 ;
        RECT 0.525 2.64 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 6.815 1.92 7.105 2.15 ;
      RECT 3.455 1.92 3.745 2.15 ;
      RECT 1.055 1.92 1.345 2.15 ;
      RECT 1.055 1.965 7.105 2.105 ;
    LAYER li ;
      RECT 9.165 0.43 9.39 2.49 ;
      RECT 9.165 1.335 10.035 1.665 ;
      RECT 9.165 0.43 9.525 1.665 ;
      RECT 8.16 2.095 8.465 2.96 ;
      RECT 7.565 2.095 8.465 2.425 ;
      RECT 7.565 2.095 8.995 2.265 ;
      RECT 8.825 0.695 8.995 2.265 ;
      RECT 8.3 0.695 8.995 1.025 ;
      RECT 6.37 2.265 6.695 2.735 ;
      RECT 6.515 0.695 6.695 2.735 ;
      RECT 8.395 1.195 8.655 1.865 ;
      RECT 6.515 1.195 8.655 1.365 ;
      RECT 6.515 0.695 6.775 1.365 ;
      RECT 0.095 2.3 0.355 2.97 ;
      RECT 0.095 2.3 0.835 2.47 ;
      RECT 0.665 1.1 0.835 2.47 ;
      RECT 6.105 1.755 6.345 2.085 ;
      RECT 6.175 0.255 6.345 2.085 ;
      RECT 0.665 1.1 1.125 1.77 ;
      RECT 0.955 0.28 1.125 1.77 ;
      RECT 3.225 0.47 3.395 1.605 ;
      RECT 1.655 1.175 2.685 1.345 ;
      RECT 2.515 0.47 2.685 1.345 ;
      RECT 0.095 1.1 1.125 1.28 ;
      RECT 1.655 0.28 1.825 1.345 ;
      RECT 0.095 0.62 0.425 1.28 ;
      RECT 4.47 0.525 6.345 0.705 ;
      RECT 2.515 0.47 4.835 0.64 ;
      RECT 5.505 0.255 7.175 0.525 ;
      RECT 0.955 0.28 1.825 0.45 ;
      RECT 5.765 2.265 6.2 2.465 ;
      RECT 5.765 0.875 5.935 2.465 ;
      RECT 4.225 1.355 4.555 1.955 ;
      RECT 4.225 1.495 5.935 1.665 ;
      RECT 5.665 0.875 5.935 1.665 ;
      RECT 5.665 0.875 5.995 1.065 ;
      RECT 5.155 0.93 5.485 1.315 ;
      RECT 3.565 0.93 5.485 1.14 ;
      RECT 3.565 0.81 4.145 1.14 ;
      RECT 2.81 2.845 3.585 3.075 ;
      RECT 3.415 2.445 3.585 3.075 ;
      RECT 4.145 2.445 4.415 3.035 ;
      RECT 4.195 2.125 4.415 3.035 ;
      RECT 3.415 2.445 4.415 2.615 ;
      RECT 4.195 2.125 5.485 2.295 ;
      RECT 5.155 1.845 5.485 2.295 ;
      RECT 3.455 1.875 4.015 2.18 ;
      RECT 3.685 1.31 4.015 2.18 ;
      RECT 2.41 2.505 2.64 3.035 ;
      RECT 1.48 2.505 1.74 3.035 ;
      RECT 1.48 2.505 3.245 2.675 ;
      RECT 3.075 1.785 3.245 2.675 ;
      RECT 2.855 1.785 3.245 1.955 ;
      RECT 2.855 0.81 3.055 1.955 ;
      RECT 1.025 1.94 1.285 2.96 ;
      RECT 1.025 2.135 2.905 2.335 ;
      RECT 1.025 1.94 1.485 2.335 ;
      RECT 1.295 0.62 1.485 2.335 ;
      RECT 6.865 1.545 7.055 2.215 ;
  END
END scs130lp_dfrtp_1

MACRO scs130lp_dfrtp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfrtp_2 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.45 0.47 2.12 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 1.21 2.325 1.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.23 0.255 10.455 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.035 1.745 8.495 2.255 ;
        RECT 7.215 1.745 8.495 2.015 ;
        RECT 6.865 2.295 7.385 2.605 ;
        RECT 7.215 1.745 7.385 2.605 ;
        RECT 5.495 2.905 7.035 3.075 ;
        RECT 6.865 2.295 7.035 3.075 ;
        RECT 5.495 2.235 5.665 3.075 ;
        RECT 4.625 2.235 5.665 2.565 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 10.625 -0.085 10.92 1.095 ;
        RECT 9.705 -0.085 10.06 1.015 ;
        RECT 9.57 -0.085 10.06 0.475 ;
        RECT 7.51 -0.085 7.84 0.885 ;
        RECT 5.045 -0.085 5.315 0.635 ;
        RECT 1.995 -0.085 2.24 0.7 ;
        RECT 0.56 -0.085 0.785 0.88 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.04 3.415 ;
        RECT 10.625 1.815 10.92 3.415 ;
        RECT 9.725 1.815 10.06 3.415 ;
        RECT 8.7 2.775 9.03 3.415 ;
        RECT 7.205 2.775 8.16 3.415 ;
        RECT 5.065 2.735 5.325 3.415 ;
        RECT 3.755 2.72 3.995 3.415 ;
        RECT 1.98 2.765 2.31 3.415 ;
        RECT 0.525 2.64 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 6.815 1.55 7.105 1.78 ;
      RECT 3.455 1.55 3.745 1.78 ;
      RECT 1.535 1.55 1.825 1.78 ;
      RECT 1.535 1.595 7.105 1.735 ;
    LAYER li ;
      RECT 9.22 2.515 9.555 3.075 ;
      RECT 9.365 1.185 9.555 3.075 ;
      RECT 9.365 1.185 10.06 1.515 ;
      RECT 9.365 0.645 9.535 3.075 ;
      RECT 9.14 0.255 9.4 0.815 ;
      RECT 8.33 2.435 8.53 3.05 ;
      RECT 7.575 2.435 8.835 2.605 ;
      RECT 8.665 2.175 8.835 2.605 ;
      RECT 7.575 2.185 7.825 2.605 ;
      RECT 8.665 2.175 9.195 2.345 ;
      RECT 9.025 0.985 9.195 2.345 ;
      RECT 8.3 0.985 9.195 1.155 ;
      RECT 8.3 0.67 8.63 1.155 ;
      RECT 6.265 2.405 6.695 2.735 ;
      RECT 6.525 0.605 6.695 2.735 ;
      RECT 8.685 1.325 8.855 1.995 ;
      RECT 7.225 1.325 8.855 1.495 ;
      RECT 7.225 1.055 7.395 1.495 ;
      RECT 6.525 1.055 7.395 1.225 ;
      RECT 6.525 0.605 6.775 1.225 ;
      RECT 0.095 2.3 0.355 2.97 ;
      RECT 0.095 2.3 0.835 2.47 ;
      RECT 0.665 1.1 0.835 2.47 ;
      RECT 6.175 0.255 6.355 2.075 ;
      RECT 0.665 1.1 1.125 1.705 ;
      RECT 0.955 0.255 1.125 1.705 ;
      RECT 3.135 1.14 3.5 1.385 ;
      RECT 3.33 0.255 3.5 1.385 ;
      RECT 0.095 1.1 1.125 1.27 ;
      RECT 0.095 0.545 0.39 1.27 ;
      RECT 1.655 0.87 2.58 1.04 ;
      RECT 2.41 0.255 2.58 1.04 ;
      RECT 4.05 0.805 5.655 0.975 ;
      RECT 5.485 0.255 5.655 0.975 ;
      RECT 1.655 0.255 1.825 1.04 ;
      RECT 4.05 0.255 4.22 0.975 ;
      RECT 2.41 0.255 4.22 0.47 ;
      RECT 6.175 0.255 7.175 0.435 ;
      RECT 5.485 0.255 7.175 0.425 ;
      RECT 0.955 0.255 1.825 0.425 ;
      RECT 5.835 2.405 6.095 2.735 ;
      RECT 5.835 0.595 6.005 2.735 ;
      RECT 4.265 1.495 6.005 1.675 ;
      RECT 5.825 0.595 6.005 1.675 ;
      RECT 3.67 1.145 5.645 1.325 ;
      RECT 3.67 0.64 3.88 1.325 ;
      RECT 4.165 1.92 4.455 3.05 ;
      RECT 2.87 2.765 3.585 3.05 ;
      RECT 3.415 1.92 3.585 3.05 ;
      RECT 3.415 1.92 4.455 2.22 ;
      RECT 4.185 1.845 5.645 2.065 ;
      RECT 2.48 2.425 2.7 3.05 ;
      RECT 1.55 2.425 1.81 3.05 ;
      RECT 1.55 2.425 3.245 2.595 ;
      RECT 3.075 1.565 3.245 2.595 ;
      RECT 2.785 1.565 3.245 1.735 ;
      RECT 2.785 0.64 2.955 1.735 ;
      RECT 2.785 0.64 3.16 0.97 ;
      RECT 1.025 2.085 1.285 2.97 ;
      RECT 1.025 2.085 2.905 2.255 ;
      RECT 2.645 1.925 2.905 2.255 ;
      RECT 1.295 0.595 1.475 2.255 ;
      RECT 1.295 1.5 1.825 1.83 ;
      RECT 1.295 0.595 1.485 1.83 ;
      RECT 6.865 1.455 7.045 2.125 ;
      RECT 3.415 1.555 4.005 1.75 ;
  END
END scs130lp_dfrtp_2

MACRO scs130lp_dfrtp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfrtp_4 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.2 0.47 2.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.455 2.82 1.85 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.31 1.755 11.85 1.925 ;
        RECT 11.68 1.065 11.85 1.925 ;
        RECT 10.31 1.065 11.85 1.235 ;
        RECT 11.205 1.755 11.395 3.075 ;
        RECT 11.15 0.255 11.395 1.235 ;
        RECT 10.31 1.755 10.535 3.075 ;
        RECT 10.31 0.255 10.535 1.235 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.155 1.45 8.565 2.12 ;
        RECT 7.345 1.45 8.565 1.62 ;
        RECT 5.785 2.785 7.515 2.955 ;
        RECT 7.345 1.45 7.515 2.955 ;
        RECT 4.895 2.635 5.955 2.805 ;
        RECT 4.895 2.255 5.065 2.805 ;
        RECT 4.735 2.255 5.065 2.52 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12 0.085 ;
        RECT 11.565 -0.085 11.895 0.895 ;
        RECT 10.705 -0.085 10.98 0.895 ;
        RECT 9.88 -0.085 10.14 1.095 ;
        RECT 7.895 -0.085 8.225 0.93 ;
        RECT 5.155 -0.085 5.485 0.355 ;
        RECT 2.235 -0.085 2.48 0.915 ;
        RECT 0.525 -0.085 0.865 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
      LAYER li ;
        RECT 0 3.245 12 3.415 ;
        RECT 11.565 2.095 11.895 3.415 ;
        RECT 10.705 2.095 11.035 3.415 ;
        RECT 9.88 1.815 10.14 3.415 ;
        RECT 8.875 2.64 9.205 3.415 ;
        RECT 7.715 2.64 8.045 3.415 ;
        RECT 5.275 2.975 5.605 3.415 ;
        RECT 3.935 2.795 4.15 3.415 ;
        RECT 2.09 2.795 2.42 3.415 ;
        RECT 0.625 2.64 0.935 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 6.815 1.92 7.105 2.15 ;
      RECT 3.935 1.92 4.225 2.15 ;
      RECT 1.055 1.92 1.345 2.15 ;
      RECT 1.055 1.965 7.105 2.105 ;
    LAYER li ;
      RECT 9.465 0.255 9.71 3.075 ;
      RECT 9.465 1.405 11.5 1.585 ;
      RECT 8.365 2.3 8.695 2.815 ;
      RECT 7.685 2.3 9.295 2.47 ;
      RECT 9.125 0.65 9.295 2.47 ;
      RECT 7.685 1.95 7.945 2.47 ;
      RECT 8.84 0.65 9.295 0.93 ;
      RECT 6.33 2.345 6.66 2.615 ;
      RECT 6.485 1.595 6.66 2.615 ;
      RECT 8.735 1.1 8.955 1.865 ;
      RECT 6.655 0.865 6.845 1.765 ;
      RECT 6.655 1.1 8.955 1.27 ;
      RECT 6.655 0.865 6.985 1.27 ;
      RECT 0.195 2.3 0.455 2.97 ;
      RECT 0.195 2.3 0.935 2.47 ;
      RECT 0.765 0.86 0.935 2.47 ;
      RECT 6.125 1.245 6.315 1.955 ;
      RECT 0.765 0.86 1.205 1.65 ;
      RECT 1.035 0.29 1.205 1.65 ;
      RECT 3.365 1.235 3.59 1.565 ;
      RECT 3.42 0.365 3.59 1.565 ;
      RECT 6.315 0.525 6.485 1.415 ;
      RECT 1.895 1.085 2.82 1.255 ;
      RECT 2.65 0.365 2.82 1.255 ;
      RECT 1.895 0.29 2.065 1.255 ;
      RECT 0.095 0.86 1.205 1.03 ;
      RECT 0.095 0.495 0.355 1.03 ;
      RECT 4.14 0.525 7.425 0.695 ;
      RECT 7.095 0.255 7.425 0.695 ;
      RECT 2.65 0.365 4.31 0.535 ;
      RECT 1.035 0.29 2.065 0.46 ;
      RECT 5.785 2.205 6.15 2.465 ;
      RECT 5.785 0.865 5.955 2.465 ;
      RECT 4.375 1.215 4.705 1.745 ;
      RECT 4.375 1.485 5.955 1.655 ;
      RECT 5.785 0.865 6.145 1.065 ;
      RECT 5.275 0.875 5.605 1.315 ;
      RECT 3.76 0.875 5.605 1.045 ;
      RECT 3.76 0.715 3.96 1.045 ;
      RECT 2.99 2.795 3.765 3.075 ;
      RECT 3.595 2.455 3.765 3.075 ;
      RECT 4.32 2.625 4.585 3.05 ;
      RECT 3.595 2.455 4.545 2.625 ;
      RECT 4.375 1.915 4.545 3.05 ;
      RECT 4.375 1.915 5.605 2.085 ;
      RECT 5.275 1.825 5.605 2.085 ;
      RECT 2.59 2.455 2.82 3.05 ;
      RECT 1.66 2.455 1.92 3.05 ;
      RECT 1.66 2.455 3.425 2.625 ;
      RECT 3.255 1.745 3.425 2.625 ;
      RECT 2.99 1.745 3.425 1.915 ;
      RECT 2.99 0.725 3.195 1.915 ;
      RECT 2.99 0.725 3.25 1.055 ;
      RECT 1.105 1.87 1.385 2.96 ;
      RECT 1.105 2.085 3.085 2.285 ;
      RECT 1.385 0.63 1.715 2.285 ;
      RECT 6.83 1.935 7.165 2.195 ;
      RECT 3.835 1.215 4.205 2.18 ;
  END
END scs130lp_dfrtp_4

MACRO scs130lp_dfsbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfsbp_1 0 0 ;
  SIZE 12.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.47 2.09 ;
        RECT 0.085 1.21 0.43 2.49 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 2.175 2.55 2.505 ;
        RECT 2 1.355 2.425 2.505 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.04 0.47 11.41 2.225 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.94 1.74 12.395 3.075 ;
        RECT 12.125 0.26 12.395 3.075 ;
    END
  END QN
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.51 1.715 8.365 2.045 ;
        RECT 6.33 2.845 7.68 3.075 ;
        RECT 7.51 1.715 7.68 3.075 ;
        RECT 6.33 2.245 6.5 3.075 ;
        RECT 5.165 2.245 6.5 2.49 ;
        RECT 5.165 1.945 5.495 2.49 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.48 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.48 0.085 ;
        RECT 11.58 -0.085 11.91 1.06 ;
        RECT 9.605 -0.085 9.865 0.97 ;
        RECT 8.62 -0.085 8.95 0.73 ;
        RECT 5.25 -0.085 5.52 1.075 ;
        RECT 3.725 -0.085 3.925 0.905 ;
        RECT 1.645 -0.085 1.975 0.845 ;
        RECT 0.1 -0.085 0.43 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.48 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.48 3.415 ;
        RECT 11.44 2.735 11.77 3.415 ;
        RECT 9.57 2.155 9.885 3.415 ;
        RECT 7.85 2.28 8.09 3.415 ;
        RECT 5.82 2.66 6.15 3.415 ;
        RECT 3.77 2.825 4.1 3.415 ;
        RECT 2 2.675 2.33 3.415 ;
        RECT 0.1 2.66 0.43 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.81 2.285 7.14 2.675 ;
      RECT 6.935 1.315 7.14 2.675 ;
      RECT 10.7 2.395 11.75 2.565 ;
      RECT 11.58 1.23 11.75 2.565 ;
      RECT 8.29 2.225 8.705 2.555 ;
      RECT 8.535 1.315 8.705 2.555 ;
      RECT 10.7 1.325 10.87 2.565 ;
      RECT 9.265 1.315 9.595 1.985 ;
      RECT 11.58 1.23 11.955 1.56 ;
      RECT 9.265 1.325 10.87 1.495 ;
      RECT 6.935 1.315 9.595 1.485 ;
      RECT 6.935 0.955 7.105 2.675 ;
      RECT 6.7 0.955 7.105 1.165 ;
      RECT 10.055 1.985 10.34 2.805 ;
      RECT 10.28 1.665 10.53 2.155 ;
      RECT 7.805 0.955 9.435 1.145 ;
      RECT 9.14 0.64 9.435 1.145 ;
      RECT 8.875 2.2 9.13 3.065 ;
      RECT 8.875 2.2 9.4 2.53 ;
      RECT 6.2 0.615 6.53 1.075 ;
      RECT 6.2 0.615 8.1 0.785 ;
      RECT 7.83 0.4 8.1 0.785 ;
      RECT 5.74 0.265 6.01 1.075 ;
      RECT 5.74 0.265 7.62 0.445 ;
      RECT 0.965 2.26 1.315 3.075 ;
      RECT 0.6 2.26 1.315 2.93 ;
      RECT 0.64 0.83 0.84 2.93 ;
      RECT 3.4 1.075 3.615 2.165 ;
      RECT 6.505 1.335 6.765 2.005 ;
      RECT 6.27 1.335 6.765 1.505 ;
      RECT 0.64 1.285 1.83 1.455 ;
      RECT 1.635 1.015 1.83 1.455 ;
      RECT 4.815 1.245 6.53 1.415 ;
      RECT 0.64 0.83 0.9 1.455 ;
      RECT 3.4 1.075 4.265 1.245 ;
      RECT 4.095 0.605 4.265 1.245 ;
      RECT 4.815 0.605 4.985 1.415 ;
      RECT 3.325 0.3 3.495 1.235 ;
      RECT 1.635 1.015 2.315 1.185 ;
      RECT 2.145 0.3 2.315 1.185 ;
      RECT 4.095 0.605 4.985 0.775 ;
      RECT 2.145 0.3 3.495 0.47 ;
      RECT 3.06 2.485 3.31 3.05 ;
      RECT 3.06 2.485 3.955 2.655 ;
      RECT 3.785 1.765 3.955 2.655 ;
      RECT 4.675 1.765 4.985 2.505 ;
      RECT 3.06 1.415 3.23 3.05 ;
      RECT 5.675 1.685 6.215 2.015 ;
      RECT 3.785 1.765 4.985 1.935 ;
      RECT 4.815 1.595 5.845 1.765 ;
      RECT 2.945 0.645 3.155 1.585 ;
      RECT 4.28 2.685 5.565 3.015 ;
      RECT 4.28 2.175 4.45 3.015 ;
      RECT 4.135 2.175 4.45 2.505 ;
      RECT 3.9 1.415 4.635 1.585 ;
      RECT 4.445 0.955 4.635 1.585 ;
      RECT 2.55 2.72 2.89 3.05 ;
      RECT 2.72 1.765 2.89 3.05 ;
      RECT 2.605 0.645 2.775 1.935 ;
      RECT 2.485 0.645 2.775 0.975 ;
      RECT 1.485 1.815 1.765 2.975 ;
      RECT 1.02 1.815 1.765 2.09 ;
      RECT 1.205 0.265 1.465 0.945 ;
      RECT 0.805 0.265 1.465 0.515 ;
      RECT 10.035 0.64 10.73 1.155 ;
  END
END scs130lp_dfsbp_1

MACRO scs130lp_dfsbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfsbp_2 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.485 0.54 2.12 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.915 1.605 2.595 2.515 ;
        RECT 1.915 1.365 2.245 2.515 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.145 0.375 12.39 3.075 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.225 0.255 10.465 3.075 ;
    END
  END QN
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.43 1.765 8.345 2.095 ;
        RECT 6.435 2.905 7.62 3.075 ;
        RECT 7.43 1.765 7.62 3.075 ;
        RECT 6.435 2.205 6.605 3.075 ;
        RECT 5.315 2.205 6.605 2.49 ;
        RECT 5.315 1.845 5.505 2.49 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.96 0.085 ;
        RECT 12.56 -0.085 12.86 1.255 ;
        RECT 11.67 -0.085 11.975 1.175 ;
        RECT 10.635 -0.085 10.98 1.095 ;
        RECT 9.765 -0.085 10.055 0.895 ;
        RECT 8.72 -0.085 9.05 0.815 ;
        RECT 5.41 -0.085 5.74 0.995 ;
        RECT 3.815 -0.085 4.075 0.955 ;
        RECT 1.73 -0.085 2.06 0.845 ;
        RECT 0.185 -0.085 0.45 1.27 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.96 3.415 ;
        RECT 12.56 1.815 12.86 3.415 ;
        RECT 11.67 1.845 11.975 3.415 ;
        RECT 10.645 1.815 10.98 3.415 ;
        RECT 9.725 2.155 10.055 3.415 ;
        RECT 7.79 2.275 8.085 3.415 ;
        RECT 5.985 2.66 6.265 3.415 ;
        RECT 3.84 2.835 4.675 3.415 ;
        RECT 2.03 2.685 2.36 3.415 ;
        RECT 0.19 2.29 0.52 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 11.15 0.7 11.465 2.485 ;
      RECT 11.15 1.345 11.975 1.675 ;
      RECT 11.15 0.7 11.48 1.675 ;
      RECT 9.2 1.815 9.53 2.21 ;
      RECT 9.2 1.815 10.005 1.985 ;
      RECT 9.835 1.065 10.005 1.985 ;
      RECT 8.025 1.065 10.005 1.235 ;
      RECT 8.025 0.985 9.57 1.235 ;
      RECT 9.24 0.7 9.57 1.235 ;
      RECT 6.785 2.405 7.25 2.735 ;
      RECT 7.08 0.975 7.25 2.735 ;
      RECT 8.255 2.275 8.695 2.605 ;
      RECT 8.525 1.405 8.695 2.605 ;
      RECT 8.525 1.405 9.655 1.645 ;
      RECT 7.08 1.405 9.655 1.585 ;
      RECT 6.835 0.975 7.25 1.175 ;
      RECT 6.365 0.635 6.665 1.17 ;
      RECT 6.365 0.635 8.26 0.805 ;
      RECT 7.93 0.5 8.26 0.805 ;
      RECT 5.91 0.265 6.17 0.995 ;
      RECT 5.91 0.265 7.74 0.465 ;
      RECT 0.72 2.775 1.215 3.075 ;
      RECT 0.72 1.015 0.95 3.075 ;
      RECT 0.69 2.29 0.95 2.63 ;
      RECT 3.465 1.125 3.655 2.185 ;
      RECT 6.65 1.355 6.91 2.025 ;
      RECT 6.025 1.355 6.91 1.525 ;
      RECT 0.72 1.015 1.675 1.485 ;
      RECT 6.025 1.165 6.195 1.525 ;
      RECT 4.975 1.165 6.195 1.335 ;
      RECT 0.62 1.015 1.675 1.305 ;
      RECT 3.465 1.125 4.425 1.295 ;
      RECT 4.255 0.515 4.425 1.295 ;
      RECT 0.62 1.015 2.41 1.195 ;
      RECT 2.24 0.255 2.41 1.195 ;
      RECT 4.975 0.515 5.145 1.335 ;
      RECT 3.465 0.255 3.645 2.185 ;
      RECT 4.255 0.515 5.145 0.72 ;
      RECT 2.24 0.255 3.645 0.425 ;
      RECT 3.115 2.365 3.375 3.045 ;
      RECT 3.115 2.365 3.995 2.535 ;
      RECT 3.825 1.815 3.995 2.535 ;
      RECT 3.115 0.67 3.295 3.045 ;
      RECT 4.65 1.815 5.145 2.325 ;
      RECT 4.975 1.505 5.145 2.325 ;
      RECT 5.675 1.705 6.41 2.035 ;
      RECT 3.825 1.815 5.145 1.985 ;
      RECT 5.675 1.505 5.845 2.035 ;
      RECT 4.975 1.505 5.845 1.675 ;
      RECT 2.985 0.67 3.295 1 ;
      RECT 4.845 2.72 5.73 3.075 ;
      RECT 4.845 2.495 5.145 3.075 ;
      RECT 4.175 2.495 5.145 2.665 ;
      RECT 4.175 2.185 4.345 2.665 ;
      RECT 3.965 1.465 4.795 1.645 ;
      RECT 4.595 0.89 4.795 1.645 ;
      RECT 2.64 2.695 2.945 3.025 ;
      RECT 2.765 1.265 2.945 3.025 ;
      RECT 2.58 0.67 2.815 1.435 ;
      RECT 1.48 2.305 1.745 2.975 ;
      RECT 1.215 1.805 1.545 2.475 ;
      RECT 0.955 0.255 1.55 0.845 ;
  END
END scs130lp_dfsbp_2

MACRO scs130lp_dfsbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfsbp_lp 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.45 1.89 1.78 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.55 1.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.215 1.85 13.805 2.89 ;
        RECT 13.635 0.265 13.805 2.89 ;
        RECT 13.475 0.265 13.805 0.725 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.595 1.18 11.925 3.02 ;
        RECT 11.495 0.265 11.665 1.78 ;
        RECT 11.335 0.265 11.665 0.725 ;
    END
  END QN
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
      ANTENNAGATEAREA 0.626 LAYER met1 ;
      ANTENNAMAXAREACAR 1.046166 LAYER li ;
      ANTENNAMAXAREACAR 1.046166 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.801917 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.801917 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.092332 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 9.695 1.92 9.985 2.15 ;
        RECT 6.335 1.965 9.985 2.105 ;
        RECT 6.335 1.92 6.625 2.15 ;
      LAYER li ;
        RECT 9.585 1.265 9.955 2.15 ;
        RECT 6.395 1.605 6.665 2.15 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.92 0.085 ;
        RECT 12.685 -0.085 13.015 0.725 ;
        RECT 10.545 -0.085 10.875 0.725 ;
        RECT 8.945 -0.085 9.275 0.735 ;
        RECT 6.75 -0.085 7.08 1.065 ;
        RECT 4.915 -0.085 5.165 0.685 ;
        RECT 2.28 -0.085 2.45 0.92 ;
        RECT 0.095 -0.085 0.425 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.92 3.415 ;
        RECT 12.685 1.85 13.015 3.415 ;
        RECT 11.145 2.02 11.395 3.415 ;
        RECT 9.11 2.68 9.44 3.415 ;
        RECT 6.495 2.855 6.825 3.415 ;
        RECT 4.985 2.855 5.315 3.415 ;
        RECT 1.825 2.31 2.155 3.415 ;
        RECT 0.17 2.025 0.5 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 12.105 1.49 12.485 2.89 ;
      RECT 12.105 1.49 13.32 1.66 ;
      RECT 12.99 0.99 13.32 1.66 ;
      RECT 12.105 0.265 12.275 2.89 ;
      RECT 11.895 0.265 12.275 0.725 ;
      RECT 9.81 2.895 10.965 3.065 ;
      RECT 10.795 1.17 10.965 3.065 ;
      RECT 7.805 2.075 8.135 3.065 ;
      RECT 9.81 2.33 10.14 3.065 ;
      RECT 7.805 2.33 10.14 2.5 ;
      RECT 8.76 0.915 8.93 2.5 ;
      RECT 10.795 1.17 11.125 1.84 ;
      RECT 7.925 0.915 8.93 1.085 ;
      RECT 7.65 0.605 8.095 1.065 ;
      RECT 10.365 0.915 10.615 2.715 ;
      RECT 9.11 0.915 9.375 1.885 ;
      RECT 9.11 0.915 10.615 1.085 ;
      RECT 9.755 0.265 10.085 1.085 ;
      RECT 2.355 2.895 4.545 3.065 ;
      RECT 4.375 2.505 4.545 3.065 ;
      RECT 3.515 1.33 3.685 3.065 ;
      RECT 2.355 2.31 2.685 3.065 ;
      RECT 4.375 2.505 7.585 2.675 ;
      RECT 7.415 1.3 7.585 2.675 ;
      RECT 8.315 1.46 8.58 1.935 ;
      RECT 2.99 1.33 4.52 1.78 ;
      RECT 7.415 1.46 8.58 1.63 ;
      RECT 7.415 1.3 7.745 1.63 ;
      RECT 2.99 0.615 3.32 1.78 ;
      RECT 3.865 2.075 4.195 2.715 ;
      RECT 3.865 2.075 4.87 2.245 ;
      RECT 4.7 0.865 4.87 2.245 ;
      RECT 6.875 1.245 7.205 1.915 ;
      RECT 5.62 1.565 6.215 1.895 ;
      RECT 6.045 1.245 6.215 1.895 ;
      RECT 6.045 1.245 7.205 1.415 ;
      RECT 6.3 0.265 6.47 1.415 ;
      RECT 4.085 0.865 4.87 1.065 ;
      RECT 4.085 0.865 5.515 1.035 ;
      RECT 5.345 0.265 5.515 1.035 ;
      RECT 4.085 0.425 4.335 1.065 ;
      RECT 5.345 0.265 6.47 0.435 ;
      RECT 5.05 2.075 6.215 2.325 ;
      RECT 5.05 1.215 5.38 2.325 ;
      RECT 5.05 1.215 5.865 1.385 ;
      RECT 5.695 0.615 5.865 1.385 ;
      RECT 5.695 0.615 6.12 1.065 ;
      RECT 0.7 2.025 1.03 3.065 ;
      RECT 0.86 0.265 1.03 3.065 ;
      RECT 3.005 1.96 3.335 2.715 ;
      RECT 2.64 1.96 3.335 2.13 ;
      RECT 2.64 0.265 2.81 2.13 ;
      RECT 1.92 1.1 2.81 1.27 ;
      RECT 1.92 0.265 2.09 1.27 ;
      RECT 3.51 0.265 3.84 0.885 ;
      RECT 0.86 0.265 1.215 0.725 ;
      RECT 2.64 0.265 3.84 0.435 ;
      RECT 0.86 0.265 2.09 0.435 ;
      RECT 1.21 1.96 1.625 3.065 ;
      RECT 1.21 1.96 2.46 2.13 ;
      RECT 2.13 1.555 2.46 2.13 ;
      RECT 1.21 0.905 1.38 3.065 ;
      RECT 1.21 0.905 1.74 1.075 ;
      RECT 1.41 0.615 1.74 1.075 ;
  END
END scs130lp_dfsbp_lp

MACRO scs130lp_dfstp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfstp_1 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 0.84 0.875 1.39 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.435 1.855 1.835 2.19 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.205 0.255 10.475 3.075 ;
        RECT 10.095 0.255 10.475 1.095 ;
    END
  END Q
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.885 1.245 7.605 1.915 ;
        RECT 4.09 1.765 6.055 1.935 ;
        RECT 4.27 0.845 4.805 1.095 ;
        RECT 4.27 0.845 4.44 1.935 ;
        RECT 4.09 1.765 4.3 2.155 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.57 -0.085 9.925 1.095 ;
        RECT 7.13 -0.085 7.46 0.735 ;
        RECT 5.065 -0.085 5.425 0.885 ;
        RECT 4.6 -0.085 5.425 0.61 ;
        RECT 3.29 -0.085 3.62 0.765 ;
        RECT 1.545 -0.085 1.845 0.97 ;
        RECT 0.665 -0.085 0.865 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.56 1.825 10.035 3.415 ;
        RECT 8.31 1.585 8.48 3.415 ;
        RECT 8.23 1.585 8.48 1.925 ;
        RECT 7.53 2.435 7.7 3.415 ;
        RECT 4.285 2.355 4.73 3.415 ;
        RECT 4.47 2.105 4.73 3.415 ;
        RECT 3.295 2.36 3.58 3.415 ;
        RECT 1.595 2.36 1.895 3.415 ;
        RECT 0.565 2.305 0.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 5.375 1.18 5.665 1.41 ;
      RECT 1.055 1.18 1.345 1.41 ;
      RECT 1.055 1.225 5.665 1.365 ;
    LAYER li ;
      RECT 9.12 0.7 9.39 2.485 ;
      RECT 9.12 1.315 10.035 1.645 ;
      RECT 8.65 0.315 8.93 3.065 ;
      RECT 7.66 0.315 7.99 0.735 ;
      RECT 7.66 0.315 8.93 0.485 ;
      RECT 7.88 2.095 8.14 2.69 ;
      RECT 5.92 2.105 6.405 2.325 ;
      RECT 7.775 0.905 8.05 2.265 ;
      RECT 6.235 2.095 8.14 2.265 ;
      RECT 7.775 0.905 8.475 1.335 ;
      RECT 8.16 0.665 8.475 1.335 ;
      RECT 5.885 0.905 8.475 1.075 ;
      RECT 5.885 0.285 6.305 1.075 ;
      RECT 5.42 2.495 7.35 2.665 ;
      RECT 7.02 2.435 7.35 2.665 ;
      RECT 5.42 2.125 5.75 2.665 ;
      RECT 4.9 2.835 6.8 3.075 ;
      RECT 4.9 2.105 5.23 3.075 ;
      RECT 5.375 1.38 5.705 1.595 ;
      RECT 5.435 1.21 5.705 1.595 ;
      RECT 3.75 2.36 4.115 2.69 ;
      RECT 3.75 1.895 3.92 2.69 ;
      RECT 3.12 1.895 3.92 2.155 ;
      RECT 3.105 0.935 3.435 1.385 ;
      RECT 3.105 0.935 4.08 1.105 ;
      RECT 3.81 0.28 4.08 1.105 ;
      RECT 2.455 2.355 2.925 2.685 ;
      RECT 2.755 0.645 2.925 2.685 ;
      RECT 2.755 1.555 3.92 1.725 ;
      RECT 3.66 1.285 3.92 1.725 ;
      RECT 2.405 0.645 2.925 0.975 ;
      RECT 2.065 2.015 2.285 2.69 ;
      RECT 2.065 2.015 2.575 2.185 ;
      RECT 2.405 1.175 2.575 2.185 ;
      RECT 2.015 1.175 2.575 1.345 ;
      RECT 2.015 0.64 2.235 1.345 ;
      RECT 1.045 0.41 1.255 2.965 ;
      RECT 2.005 1.515 2.235 1.845 ;
      RECT 1.045 1.515 2.235 1.685 ;
      RECT 1.045 0.41 1.355 1.685 ;
      RECT 0.09 1.56 0.395 2.965 ;
      RECT 0.09 1.56 0.865 1.81 ;
      RECT 0.09 0.39 0.26 2.965 ;
      RECT 0.09 0.39 0.495 0.67 ;
  END
END scs130lp_dfstp_1

MACRO scs130lp_dfstp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfstp_2 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.43 0.925 0.855 1.405 ;
        RECT 0.545 0.84 0.855 1.405 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.365 1.805 1.775 2.19 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.225 0.255 10.465 3.075 ;
    END
  END Q
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.905 1.245 7.635 1.915 ;
        RECT 3.975 1.895 6.085 1.935 ;
        RECT 4.135 1.765 7.635 1.915 ;
        RECT 4.135 0.985 4.825 1.235 ;
        RECT 3.975 1.895 4.305 2.155 ;
        RECT 4.135 0.985 4.305 2.155 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 10.635 -0.085 10.935 1.095 ;
        RECT 9.745 -0.085 10.055 1.015 ;
        RECT 9.685 -0.085 10.055 0.545 ;
        RECT 7.03 -0.085 7.36 0.665 ;
        RECT 4.895 -0.085 5.225 0.815 ;
        RECT 3.195 -0.085 3.525 0.845 ;
        RECT 1.545 -0.085 1.84 0.97 ;
        RECT 0.575 -0.085 0.905 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.04 3.415 ;
        RECT 10.635 1.815 10.935 3.415 ;
        RECT 9.725 1.975 9.935 3.415 ;
        RECT 8.365 1.67 8.565 3.415 ;
        RECT 7.555 2.435 7.785 3.415 ;
        RECT 4.165 2.36 4.745 3.415 ;
        RECT 4.485 2.105 4.745 3.415 ;
        RECT 3.195 2.36 3.465 3.415 ;
        RECT 1.545 2.36 1.875 3.415 ;
        RECT 0.585 2.315 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 5.375 1.18 5.665 1.41 ;
      RECT 1.055 1.18 1.345 1.41 ;
      RECT 1.055 1.225 5.665 1.365 ;
    LAYER li ;
      RECT 9.235 0.255 9.505 2.635 ;
      RECT 9.235 1.185 10.055 1.515 ;
      RECT 9.235 0.255 9.515 1.515 ;
      RECT 8.735 0.445 9.065 3.075 ;
      RECT 7.625 0.445 7.955 0.695 ;
      RECT 7.625 0.445 9.065 0.615 ;
      RECT 7.955 2.095 8.195 2.69 ;
      RECT 7.975 0.865 8.195 2.69 ;
      RECT 5.925 2.105 6.35 2.345 ;
      RECT 6.255 2.095 8.195 2.265 ;
      RECT 7.975 0.865 8.535 1.465 ;
      RECT 8.285 0.795 8.535 1.465 ;
      RECT 5.785 0.865 8.535 1.035 ;
      RECT 5.785 0.255 6.115 1.035 ;
      RECT 5.435 2.515 7.385 2.685 ;
      RECT 7.055 2.435 7.385 2.685 ;
      RECT 5.435 2.17 5.71 2.685 ;
      RECT 4.915 2.855 6.835 3.055 ;
      RECT 4.915 2.105 5.245 3.055 ;
      RECT 3.07 1.015 3.4 1.385 ;
      RECT 3.07 1.015 3.955 1.185 ;
      RECT 3.785 0.28 3.955 1.185 ;
      RECT 3.785 0.28 4.1 0.61 ;
      RECT 3.635 2.36 3.995 2.69 ;
      RECT 3.635 1.895 3.805 2.69 ;
      RECT 3.07 1.895 3.805 2.155 ;
      RECT 2.405 2.435 2.815 2.71 ;
      RECT 2.645 0.615 2.815 2.71 ;
      RECT 2.645 1.555 3.945 1.725 ;
      RECT 3.615 1.355 3.945 1.725 ;
      RECT 2.405 0.615 2.815 0.835 ;
      RECT 2.045 2.095 2.235 2.69 ;
      RECT 2.045 2.095 2.465 2.265 ;
      RECT 2.295 1.005 2.465 2.265 ;
      RECT 2.01 1.005 2.465 1.175 ;
      RECT 2.01 0.64 2.235 1.175 ;
      RECT 1.025 2.315 1.235 2.985 ;
      RECT 1.025 0.84 1.195 2.985 ;
      RECT 1.945 1.455 2.125 1.845 ;
      RECT 1.025 1.455 2.125 1.635 ;
      RECT 1.075 0.415 1.355 1.635 ;
      RECT 0.09 1.575 0.365 2.975 ;
      RECT 0.09 1.575 0.845 1.825 ;
      RECT 0.09 0.41 0.26 2.975 ;
      RECT 0.09 0.41 0.405 0.74 ;
      RECT 5.405 1.205 5.735 1.595 ;
  END
END scs130lp_dfstp_2

MACRO scs130lp_dfstp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfstp_4 0 0 ;
  SIZE 12.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.53 0.38 0.815 2.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.77 1.915 2.34 2.245 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.8 1.765 12.39 1.935 ;
        RECT 12.145 1.075 12.39 1.935 ;
        RECT 10.8 1.075 12.39 1.245 ;
        RECT 11.695 1.765 11.885 3.075 ;
        RECT 11.695 0.255 11.885 1.245 ;
        RECT 10.8 1.765 11.025 3.075 ;
        RECT 10.8 0.255 11.025 1.245 ;
    END
  END Q
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.18 1.325 8.485 1.835 ;
        RECT 4.645 1.765 6.35 1.935 ;
        RECT 4.645 0.78 5.11 1.935 ;
        RECT 4.645 0.78 4.845 2.155 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.48 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.48 0.085 ;
        RECT 12.055 -0.085 12.385 0.905 ;
        RECT 11.195 -0.085 11.525 0.905 ;
        RECT 10.37 -0.085 10.63 1.105 ;
        RECT 7.475 -0.085 8.145 0.785 ;
        RECT 5.42 -0.085 5.75 0.885 ;
        RECT 4.905 -0.085 5.75 0.61 ;
        RECT 3.575 -0.085 3.905 0.815 ;
        RECT 1.985 -0.085 2.225 0.97 ;
        RECT 0.985 -0.085 1.205 0.87 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.48 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.48 3.415 ;
        RECT 12.055 2.105 12.385 3.415 ;
        RECT 11.195 2.105 11.525 3.415 ;
        RECT 10.375 1.795 10.63 3.415 ;
        RECT 9.005 1.72 9.265 3.415 ;
        RECT 7.995 2.355 8.325 3.415 ;
        RECT 5.015 2.105 5.275 3.415 ;
        RECT 3.805 2.36 4.135 3.415 ;
        RECT 2.135 2.415 2.465 3.415 ;
        RECT 0.695 2.64 1.025 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 5.375 1.18 5.665 1.41 ;
      RECT 1.535 1.18 1.825 1.41 ;
      RECT 1.535 1.225 5.665 1.365 ;
    LAYER li ;
      RECT 9.945 1.425 10.205 3.075 ;
      RECT 9.945 1.425 11.975 1.595 ;
      RECT 9.945 0.255 10.2 3.075 ;
      RECT 9.435 0.265 9.775 3.075 ;
      RECT 8.315 0.265 8.575 0.785 ;
      RECT 8.315 0.265 9.775 0.435 ;
      RECT 8.495 2.015 8.835 2.66 ;
      RECT 8.655 0.955 8.835 2.66 ;
      RECT 6.52 2.015 6.795 2.355 ;
      RECT 6.52 2.015 8.835 2.185 ;
      RECT 8.655 0.955 9.265 1.205 ;
      RECT 8.935 0.605 9.265 1.205 ;
      RECT 6.21 0.955 9.265 1.125 ;
      RECT 6.21 0.255 6.705 1.125 ;
      RECT 5.965 2.525 7.825 2.695 ;
      RECT 7.565 2.355 7.825 2.695 ;
      RECT 5.965 2.105 6.295 2.695 ;
      RECT 5.445 2.865 7.345 3.065 ;
      RECT 5.445 2.105 5.775 3.065 ;
      RECT 4.305 2.325 4.66 2.69 ;
      RECT 4.305 1.895 4.475 2.69 ;
      RECT 3.66 1.895 4.475 2.155 ;
      RECT 3.035 2.295 3.3 2.69 ;
      RECT 3.13 0.585 3.3 2.69 ;
      RECT 3.13 1.555 4.465 1.725 ;
      RECT 4.135 1.325 4.465 1.725 ;
      RECT 2.82 0.585 3.3 0.915 ;
      RECT 3.48 0.985 3.81 1.385 ;
      RECT 3.48 0.985 4.445 1.155 ;
      RECT 4.115 0.285 4.445 1.155 ;
      RECT 2.635 1.915 2.865 2.69 ;
      RECT 2.78 1.085 2.95 2.085 ;
      RECT 2.395 1.085 2.95 1.255 ;
      RECT 2.395 0.64 2.65 1.255 ;
      RECT 1.195 2.64 1.6 2.97 ;
      RECT 1.43 0.54 1.6 2.97 ;
      RECT 1.43 1.485 2.6 1.745 ;
      RECT 1.43 0.54 1.815 1.745 ;
      RECT 1.375 0.54 1.815 0.935 ;
      RECT 0.17 2.3 0.525 2.975 ;
      RECT 0.17 2.3 1.26 2.47 ;
      RECT 1 1.495 1.26 2.47 ;
      RECT 0.17 0.54 0.36 2.975 ;
      RECT 5.37 1.15 6.01 1.595 ;
  END
END scs130lp_dfstp_4

MACRO scs130lp_dfstp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfstp_lp 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.51 1.45 1.84 1.78 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.55 1.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.805 1.85 13.325 2.89 ;
        RECT 13.085 0.35 13.325 2.89 ;
        RECT 12.995 0.35 13.325 0.81 ;
    END
  END Q
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
      ANTENNAGATEAREA 0.626 LAYER met1 ;
      ANTENNAMAXAREACAR 0.347923 LAYER li ;
      ANTENNAMAXAREACAR 0.347923 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.421725 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.421725 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.092332 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 9.695 1.55 9.985 1.78 ;
        RECT 6.335 1.595 9.985 1.735 ;
        RECT 6.335 1.55 6.625 1.78 ;
      LAYER li ;
        RECT 9.7 1.51 10.03 1.84 ;
        RECT 6.395 1.55 6.7 1.88 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.44 0.085 ;
        RECT 12.205 -0.085 12.535 0.81 ;
        RECT 10.855 -0.085 11.185 0.645 ;
        RECT 9.435 -0.085 9.765 0.98 ;
        RECT 6.685 -0.085 7.015 1.02 ;
        RECT 4.915 -0.085 5.165 0.695 ;
        RECT 2.28 -0.085 2.45 0.92 ;
        RECT 0.095 -0.085 0.425 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.44 3.415 ;
        RECT 12.275 1.85 12.605 3.415 ;
        RECT 11.265 1.675 11.515 3.415 ;
        RECT 9.145 2.37 9.475 3.415 ;
        RECT 6.685 2.41 7.015 3.415 ;
        RECT 4.94 2.785 5.27 3.415 ;
        RECT 1.84 2.31 2.17 3.415 ;
        RECT 0.12 2.025 0.45 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 11.695 1.49 12.075 2.89 ;
      RECT 11.695 1.49 12.84 1.66 ;
      RECT 12.51 0.99 12.84 1.66 ;
      RECT 11.695 0.35 11.865 2.89 ;
      RECT 11.415 0.35 11.865 0.81 ;
      RECT 9.925 2.895 11.085 3.065 ;
      RECT 10.915 0.825 11.085 3.065 ;
      RECT 8.045 2.02 8.375 3.065 ;
      RECT 9.925 2.02 10.255 3.065 ;
      RECT 8.045 2.02 10.255 2.19 ;
      RECT 8.835 0.895 9.005 2.19 ;
      RECT 10.835 0.825 11.165 1.495 ;
      RECT 7.96 0.895 9.005 1.065 ;
      RECT 7.96 0.605 8.29 1.065 ;
      RECT 10.485 1.675 10.735 2.715 ;
      RECT 9.185 1.16 9.49 1.84 ;
      RECT 10.485 1.16 10.655 2.715 ;
      RECT 9.185 1.16 10.655 1.33 ;
      RECT 10.065 0.265 10.395 1.33 ;
      RECT 5.45 2.895 6.505 3.065 ;
      RECT 6.335 2.06 6.505 3.065 ;
      RECT 2.37 2.895 4.76 3.065 ;
      RECT 4.59 2.435 4.76 3.065 ;
      RECT 5.45 2.435 5.62 3.065 ;
      RECT 3.5 1.245 3.67 3.065 ;
      RECT 2.37 2.025 2.62 3.065 ;
      RECT 4.59 2.435 5.62 2.605 ;
      RECT 6.335 2.06 7.78 2.23 ;
      RECT 7.45 1.3 7.78 2.23 ;
      RECT 7.45 1.51 8.655 1.84 ;
      RECT 3.15 1.245 3.67 1.84 ;
      RECT 3.15 1.245 4.505 1.575 ;
      RECT 3.15 0.615 3.32 1.84 ;
      RECT 2.99 0.615 3.32 0.985 ;
      RECT 3.85 2.075 4.18 2.715 ;
      RECT 3.85 2.075 4.855 2.245 ;
      RECT 4.685 0.875 4.855 2.245 ;
      RECT 5.575 1.575 5.905 1.905 ;
      RECT 6.91 1.2 7.24 1.87 ;
      RECT 5.575 1.575 6.215 1.745 ;
      RECT 6.045 1.2 6.215 1.745 ;
      RECT 6.045 1.2 7.24 1.37 ;
      RECT 6.335 0.265 6.505 1.37 ;
      RECT 4.085 0.875 4.855 1.065 ;
      RECT 4.085 0.875 5.515 1.045 ;
      RECT 5.345 0.265 5.515 1.045 ;
      RECT 4.085 0.605 4.335 1.065 ;
      RECT 5.345 0.265 6.505 0.435 ;
      RECT 5.825 2.085 6.155 2.715 ;
      RECT 5.035 2.085 6.155 2.255 ;
      RECT 5.035 1.225 5.365 2.255 ;
      RECT 5.035 1.225 5.865 1.395 ;
      RECT 5.695 0.615 5.865 1.395 ;
      RECT 5.695 0.615 6.155 1.02 ;
      RECT 0.65 2.025 0.98 3.065 ;
      RECT 0.81 0.265 0.98 3.065 ;
      RECT 2.8 2.075 3.32 2.715 ;
      RECT 2.8 1.165 2.97 2.715 ;
      RECT 2.1 1.165 2.97 1.335 ;
      RECT 2.63 0.265 2.8 1.335 ;
      RECT 1.93 0.265 2.1 1.27 ;
      RECT 1.93 1.1 2.8 1.27 ;
      RECT 3.51 0.265 3.84 1.065 ;
      RECT 0.81 0.265 1.215 0.725 ;
      RECT 2.63 0.265 3.84 0.435 ;
      RECT 0.81 0.265 2.1 0.435 ;
      RECT 1.16 1.96 1.64 3.065 ;
      RECT 1.16 1.96 2.19 2.13 ;
      RECT 2.02 1.515 2.19 2.13 ;
      RECT 1.16 1.1 1.33 3.065 ;
      RECT 2.02 1.515 2.475 1.845 ;
      RECT 1.16 1.1 1.74 1.27 ;
      RECT 1.41 0.615 1.74 1.27 ;
  END
END scs130lp_dfstp_lp

MACRO scs130lp_dfxbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfxbp_1 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.425 2.15 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.59 1.21 2.075 2.145 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.235 0.375 9.505 3.075 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.355 8.545 2.205 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 8.745 -0.085 9.015 1.255 ;
        RECT 7.775 -0.085 8.085 1.23 ;
        RECT 6.05 -0.085 6.38 0.955 ;
        RECT 3.61 -0.085 4.335 0.915 ;
        RECT 1.755 -0.085 2.075 0.975 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 8.805 2.785 9.015 3.415 ;
        RECT 7.785 2.715 8.115 3.415 ;
        RECT 6.08 1.975 6.41 3.415 ;
        RECT 3.945 2.765 4.275 3.415 ;
        RECT 1.495 2.655 1.735 3.415 ;
        RECT 0.095 2.32 0.39 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.58 1.635 6.875 2.755 ;
      RECT 6.58 2.375 9.05 2.545 ;
      RECT 8.72 1.425 9.05 2.545 ;
      RECT 6.865 0.775 7.035 2.545 ;
      RECT 5.895 1.635 7.035 1.805 ;
      RECT 6.865 1.32 7.265 1.65 ;
      RECT 5.895 1.485 6.225 1.805 ;
      RECT 6.55 0.355 6.89 0.955 ;
      RECT 7.26 1.875 7.605 2.205 ;
      RECT 7.435 0.83 7.605 2.205 ;
      RECT 7.215 0.83 7.605 1.04 ;
      RECT 7.215 0.265 7.385 1.04 ;
      RECT 7.06 0.265 7.385 0.595 ;
      RECT 5.205 1.875 5.465 2.75 ;
      RECT 5.265 1.125 5.465 2.75 ;
      RECT 6.435 1.125 6.685 1.455 ;
      RECT 5.265 1.125 6.685 1.295 ;
      RECT 5.265 0.64 5.435 2.75 ;
      RECT 5.01 0.64 5.435 0.995 ;
      RECT 1.905 2.865 3.3 3.075 ;
      RECT 3.13 1.895 3.3 3.075 ;
      RECT 1.045 2.295 1.325 2.965 ;
      RECT 1.905 2.315 2.075 3.075 ;
      RECT 3.13 2.415 5.035 2.585 ;
      RECT 4.865 1.225 5.035 2.585 ;
      RECT 1.045 2.315 2.075 2.485 ;
      RECT 1.21 0.64 1.42 2.485 ;
      RECT 2.945 1.895 3.3 2.155 ;
      RECT 4.865 1.225 5.095 1.555 ;
      RECT 3.545 1.085 3.875 1.385 ;
      RECT 3.545 1.085 4.695 1.255 ;
      RECT 4.505 0.585 4.695 1.255 ;
      RECT 2.605 2.365 2.96 2.695 ;
      RECT 2.605 1.555 2.775 2.695 ;
      RECT 2.605 1.555 4.46 1.725 ;
      RECT 4.13 1.425 4.46 1.725 ;
      RECT 2.865 0.635 3.16 1.725 ;
      RECT 2.245 0.635 2.435 2.695 ;
      RECT 2.245 0.635 2.695 0.965 ;
      RECT 0.56 2.32 0.795 2.99 ;
      RECT 0.595 0.45 0.795 2.99 ;
      RECT 0.595 1.215 1.04 1.885 ;
      RECT 0.595 0.45 0.875 1.885 ;
      RECT 3.495 1.895 4.695 2.235 ;
  END
END scs130lp_dfxbp_1

MACRO scs130lp_dfxbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfxbp_2 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 0.84 0.47 1.795 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 1.125 2.255 2.12 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.735 0.255 9.955 3.075 ;
        RECT 9.72 0.255 9.955 1.14 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.64 0.885 8.97 3.075 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 10.125 -0.085 10.42 1.125 ;
        RECT 9.15 -0.085 9.48 0.375 ;
        RECT 8.095 -0.085 8.425 0.375 ;
        RECT 5.97 -0.085 6.49 0.975 ;
        RECT 3.475 -0.085 4.355 0.835 ;
        RECT 1.645 -0.085 1.975 0.955 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 10.125 1.815 10.415 3.415 ;
        RECT 9.15 1.82 9.48 3.415 ;
        RECT 8.045 1.815 8.47 3.415 ;
        RECT 6.27 2.335 6.73 3.415 ;
        RECT 3.945 2.575 4.275 3.415 ;
        RECT 1.58 2.64 1.83 3.415 ;
        RECT 0.095 2.28 0.405 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.9 1.985 7.17 3.075 ;
      RECT 6.965 1.255 7.17 3.075 ;
      RECT 5.995 1.985 7.17 2.165 ;
      RECT 5.995 1.505 6.325 2.165 ;
      RECT 9.37 1.32 9.555 1.65 ;
      RECT 6.965 1.255 7.435 1.515 ;
      RECT 9.37 0.545 9.54 1.65 ;
      RECT 6.965 0.355 7.135 3.075 ;
      RECT 6.66 0.355 7.135 0.975 ;
      RECT 6.66 0.545 9.54 0.715 ;
      RECT 7.545 1.83 7.875 2.485 ;
      RECT 7.545 1.815 7.815 2.485 ;
      RECT 7.605 0.895 7.815 2.485 ;
      RECT 7.605 0.895 8.47 1.625 ;
      RECT 7.545 0.895 8.47 1.085 ;
      RECT 5.315 0.64 5.565 2.705 ;
      RECT 6.535 1.145 6.795 1.815 ;
      RECT 5.315 1.145 6.795 1.315 ;
      RECT 5.075 0.64 5.565 0.975 ;
      RECT 2 2.905 3.475 3.075 ;
      RECT 3.305 1.895 3.475 3.075 ;
      RECT 1.14 2.295 1.41 2.965 ;
      RECT 2 2.3 2.17 3.075 ;
      RECT 1.14 2.3 2.17 2.47 ;
      RECT 3.305 2.235 5.145 2.405 ;
      RECT 4.955 1.175 5.145 2.405 ;
      RECT 1.215 0.64 1.475 2.47 ;
      RECT 3.125 1.895 3.475 2.155 ;
      RECT 4.455 1.005 4.785 2.065 ;
      RECT 4.525 0.585 4.785 2.065 ;
      RECT 3.485 1.005 3.815 1.385 ;
      RECT 3.485 1.005 4.785 1.175 ;
      RECT 2.765 2.405 3.125 2.735 ;
      RECT 2.765 0.64 2.945 2.735 ;
      RECT 2.765 1.555 4.285 1.725 ;
      RECT 4.025 1.355 4.285 1.725 ;
      RECT 2.765 0.64 3.015 1.725 ;
      RECT 2.35 2.3 2.595 2.63 ;
      RECT 2.425 0.625 2.595 2.63 ;
      RECT 2.18 0.625 2.595 0.955 ;
      RECT 0.575 1.93 0.855 2.95 ;
      RECT 0.79 0.33 1.04 2.1 ;
      RECT 0.595 0.33 1.04 0.72 ;
  END
END scs130lp_dfxbp_2

MACRO scs130lp_dfxbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfxbp_lp 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 0.44 0.93 1.285 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.525 1.315 1.855 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.225 0.905 9.925 1.075 ;
        RECT 9.595 0.615 9.925 1.075 ;
        RECT 9.225 0.905 9.555 2.89 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.515 0.265 12.845 3.065 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.96 0.085 ;
        RECT 11.725 -0.085 12.055 0.725 ;
        RECT 10.465 -0.085 10.715 1.075 ;
        RECT 8.335 -0.085 8.585 0.725 ;
        RECT 5.66 -0.085 5.91 1.065 ;
        RECT 3.28 -0.085 3.61 0.785 ;
        RECT 1.11 -0.085 1.36 0.865 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.96 3.415 ;
        RECT 11.985 2.115 12.315 3.415 ;
        RECT 9.755 1.815 10.085 3.415 ;
        RECT 7.795 2.37 8.125 3.415 ;
        RECT 5.49 2.465 5.82 3.415 ;
        RECT 3.865 1.985 4.195 3.415 ;
        RECT 0.64 2.775 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 10.285 1.765 10.615 2.855 ;
      RECT 10.285 1.765 12.335 1.935 ;
      RECT 12.005 1.215 12.335 1.935 ;
      RECT 12.005 0.905 12.175 1.935 ;
      RECT 11.175 0.905 12.175 1.075 ;
      RECT 11.175 0.615 11.505 1.075 ;
      RECT 8.59 2.02 9.045 3.065 ;
      RECT 8.875 0.265 9.045 3.065 ;
      RECT 7.795 2.02 9.045 2.19 ;
      RECT 7.795 1.615 8.125 2.19 ;
      RECT 9.735 1.255 11.765 1.585 ;
      RECT 10.105 0.265 10.275 1.585 ;
      RECT 8.875 0.265 9.375 0.725 ;
      RECT 8.875 0.265 10.275 0.435 ;
      RECT 6.67 2.115 7 3.065 ;
      RECT 6.67 2.115 7.615 2.285 ;
      RECT 7.445 1.265 7.615 2.285 ;
      RECT 8.365 1.17 8.695 1.84 ;
      RECT 6.92 1.265 8.695 1.435 ;
      RECT 6.92 0.965 7.09 1.435 ;
      RECT 6.14 0.265 6.39 1.155 ;
      RECT 7.825 0.265 8.155 0.725 ;
      RECT 6.14 0.265 8.155 0.435 ;
      RECT 6.14 2.075 6.47 3.065 ;
      RECT 4.395 1.755 4.78 2.755 ;
      RECT 4.61 0.965 4.78 2.755 ;
      RECT 4.395 2.115 6.47 2.285 ;
      RECT 5.31 1.335 6.74 1.505 ;
      RECT 6.57 0.615 6.74 1.505 ;
      RECT 3.075 0.965 3.405 1.455 ;
      RECT 5.31 0.265 5.48 1.505 ;
      RECT 3.075 0.965 4.78 1.135 ;
      RECT 7.27 0.615 7.6 1.085 ;
      RECT 4.15 0.265 4.48 1.135 ;
      RECT 6.57 0.615 7.6 0.785 ;
      RECT 4.15 0.265 5.48 0.435 ;
      RECT 6.935 1.615 7.265 1.935 ;
      RECT 4.96 1.685 5.29 1.935 ;
      RECT 4.96 1.685 7.265 1.855 ;
      RECT 4.96 0.615 5.13 1.935 ;
      RECT 4.71 0.615 5.13 0.785 ;
      RECT 2.25 1.595 2.58 1.855 ;
      RECT 2.25 1.635 4.215 1.805 ;
      RECT 4.045 1.315 4.215 1.805 ;
      RECT 2.33 0.405 2.66 1.805 ;
      RECT 4.045 1.315 4.43 1.575 ;
      RECT 3.335 1.985 3.665 2.755 ;
      RECT 1.72 2.425 3.665 2.595 ;
      RECT 1.72 2.385 2.05 2.595 ;
      RECT 2.78 1.985 3.11 2.245 ;
      RECT 1.17 2.035 1.5 2.245 ;
      RECT 1.17 2.035 3.11 2.205 ;
      RECT 1.82 0.405 1.99 2.205 ;
      RECT 1.82 0.405 2.15 0.865 ;
      RECT 1.15 2.775 2.315 3.065 ;
      RECT 0.11 1.995 0.44 3.035 ;
      RECT 1.15 2.425 1.32 3.065 ;
      RECT 0.11 2.425 1.32 2.595 ;
      RECT 0.11 0.405 0.42 3.035 ;
  END
END scs130lp_dfxbp_lp

MACRO scs130lp_dfxtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfxtp_1 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.425 2.155 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.58 1.21 2.075 1.79 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.775 0.255 8.065 3.075 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.34 -0.085 7.605 1.095 ;
        RECT 5.975 -0.085 6.305 0.945 ;
        RECT 3.57 -0.085 4.24 0.935 ;
        RECT 1.71 -0.085 2.04 1.04 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.305 1.825 7.605 3.415 ;
        RECT 5.98 1.965 6.36 3.415 ;
        RECT 3.76 2.635 4.09 3.415 ;
        RECT 1.51 2.3 1.735 3.415 ;
        RECT 0.095 2.325 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.54 1.625 6.935 2.75 ;
      RECT 5.79 1.625 6.935 1.795 ;
      RECT 6.765 1.27 7.605 1.655 ;
      RECT 5.79 1.465 6.12 1.795 ;
      RECT 6.765 0.945 7.17 1.655 ;
      RECT 6.475 0.415 6.935 0.945 ;
      RECT 5.11 1.875 5.375 2.755 ;
      RECT 5.205 0.64 5.375 2.755 ;
      RECT 6.335 1.125 6.595 1.455 ;
      RECT 5.205 1.125 6.595 1.295 ;
      RECT 5.205 0.64 5.395 1.295 ;
      RECT 4.99 0.64 5.395 0.97 ;
      RECT 1.905 2.605 3.495 2.88 ;
      RECT 3.325 2.285 3.495 2.88 ;
      RECT 1.045 2.045 1.34 2.715 ;
      RECT 2.595 1.575 2.775 2.88 ;
      RECT 1.905 1.96 2.075 2.88 ;
      RECT 3.325 2.285 4.93 2.455 ;
      RECT 4.76 1.425 4.93 2.455 ;
      RECT 1.18 1.96 2.075 2.13 ;
      RECT 1.18 0.855 1.41 2.13 ;
      RECT 4.855 1.195 5.035 1.595 ;
      RECT 3.37 1.855 4.58 2.115 ;
      RECT 4.41 0.575 4.58 2.115 ;
      RECT 3.37 1.445 3.7 2.115 ;
      RECT 4.41 0.575 4.685 1.245 ;
      RECT 2.945 1.105 3.155 2.435 ;
      RECT 3.98 1.105 4.24 1.675 ;
      RECT 2.945 1.105 4.24 1.275 ;
      RECT 2.755 0.86 3.125 1.19 ;
      RECT 2.245 0.86 2.425 2.435 ;
      RECT 2.245 0.86 2.575 1.19 ;
      RECT 0.595 0.4 0.795 2.99 ;
      RECT 0.595 0.955 1.01 1.625 ;
      RECT 0.595 0.4 0.855 1.625 ;
  END
END scs130lp_dfxtp_1

MACRO scs130lp_dfxtp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfxtp_2 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.425 2.49 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.94 1.14 2.27 1.765 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.785 0.375 8.05 3.075 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.64 0.085 ;
        RECT 8.22 -0.085 8.455 1.255 ;
        RECT 7.335 -0.085 7.615 1.255 ;
        RECT 6 -0.085 6.52 0.945 ;
        RECT 3.52 -0.085 4.425 0.885 ;
        RECT 1.755 -0.085 2.035 0.97 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.64 3.415 ;
        RECT 8.22 1.815 8.455 3.415 ;
        RECT 7.335 1.815 7.615 3.415 ;
        RECT 6.15 1.975 6.53 3.415 ;
        RECT 3.975 2.625 4.305 3.415 ;
        RECT 1.59 2.285 1.92 3.415 ;
        RECT 0.095 2.66 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.75 1.635 7.165 2.755 ;
      RECT 6.995 0.415 7.165 2.755 ;
      RECT 6.025 1.635 7.165 1.805 ;
      RECT 6.995 1.425 7.435 1.645 ;
      RECT 6.025 1.465 6.355 1.805 ;
      RECT 6.69 0.415 7.165 0.945 ;
      RECT 5.335 1.875 5.655 2.755 ;
      RECT 5.485 0.645 5.655 2.755 ;
      RECT 6.565 1.125 6.825 1.455 ;
      RECT 5.485 1.125 6.825 1.295 ;
      RECT 5.145 0.645 5.655 1.125 ;
      RECT 2.09 2.76 3.69 2.94 ;
      RECT 3.52 2.285 3.69 2.94 ;
      RECT 1.21 0.64 1.42 2.865 ;
      RECT 2.8 1.385 2.97 2.94 ;
      RECT 2.09 1.935 2.27 2.94 ;
      RECT 3.52 2.285 5.165 2.455 ;
      RECT 4.985 1.295 5.165 2.455 ;
      RECT 1.21 1.935 2.27 2.105 ;
      RECT 1.21 0.64 1.585 2.105 ;
      RECT 4.985 1.295 5.305 1.555 ;
      RECT 4.975 1.295 5.305 1.475 ;
      RECT 3.605 1.915 4.815 2.115 ;
      RECT 4.595 0.585 4.805 2.115 ;
      RECT 3.605 1.405 3.935 2.115 ;
      RECT 3.14 1.055 3.35 2.59 ;
      RECT 4.175 1.055 4.425 1.675 ;
      RECT 3.14 1.055 4.425 1.225 ;
      RECT 3.14 0.865 3.34 2.59 ;
      RECT 2.79 0.865 3.34 1.035 ;
      RECT 2.79 0.64 3.06 1.035 ;
      RECT 2.44 1.22 2.63 2.59 ;
      RECT 2.44 0.64 2.62 2.59 ;
      RECT 2.225 0.64 2.62 0.97 ;
      RECT 0.595 0.33 1.04 3.05 ;
  END
END scs130lp_dfxtp_2

MACRO scs130lp_dfxtp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfxtp_4 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.425 2.49 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.58 1.125 2.075 1.795 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.795 0.84 9.035 2.49 ;
        RECT 8.32 1.735 9.035 1.945 ;
        RECT 7.42 1.055 9.035 1.225 ;
        RECT 8.32 0.84 9.035 1.225 ;
        RECT 8.32 1.735 8.51 3.075 ;
        RECT 8.32 0.255 8.51 1.225 ;
        RECT 7.425 1.735 9.035 1.905 ;
        RECT 7.425 1.735 7.65 3.075 ;
        RECT 7.42 0.255 7.65 1.225 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 8.68 -0.085 9.01 0.67 ;
        RECT 7.82 -0.085 8.15 0.885 ;
        RECT 6.96 -0.085 7.25 1.095 ;
        RECT 5.785 -0.085 6.115 0.845 ;
        RECT 3.705 -0.085 4.035 0.935 ;
        RECT 1.65 -0.085 1.98 0.955 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 8.68 2.66 9.01 3.415 ;
        RECT 7.82 2.075 8.15 3.415 ;
        RECT 6.96 1.815 7.255 3.415 ;
        RECT 6.01 2.035 6.34 3.415 ;
        RECT 3.76 2.625 4.09 3.415 ;
        RECT 1.535 2.395 1.725 3.415 ;
        RECT 0.095 2.665 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.51 1.695 6.75 3.005 ;
      RECT 6.58 0.285 6.75 3.005 ;
      RECT 5.56 1.695 6.75 1.865 ;
      RECT 5.56 1.355 5.89 1.865 ;
      RECT 6.58 1.395 8.615 1.565 ;
      RECT 6.295 0.285 6.75 0.845 ;
      RECT 5.11 1.015 5.36 2.7 ;
      RECT 6.15 1.015 6.41 1.515 ;
      RECT 5.11 1.015 6.41 1.185 ;
      RECT 5.11 0.64 5.28 2.7 ;
      RECT 4.895 0.64 5.28 0.995 ;
      RECT 1.045 2.045 1.315 2.715 ;
      RECT 1.905 2.535 3.495 2.705 ;
      RECT 3.325 2.285 3.495 2.705 ;
      RECT 2.595 1.545 2.775 2.705 ;
      RECT 1.905 2.045 2.075 2.705 ;
      RECT 3.325 2.285 4.93 2.455 ;
      RECT 4.76 1.225 4.93 2.455 ;
      RECT 1.045 2.045 2.075 2.215 ;
      RECT 1.2 0.64 1.41 2.215 ;
      RECT 4.73 1.225 4.93 1.555 ;
      RECT 1.2 0.64 1.48 0.96 ;
      RECT 3.42 1.915 4.58 2.115 ;
      RECT 3.42 1.855 4.56 2.115 ;
      RECT 4.39 0.585 4.56 2.115 ;
      RECT 3.42 1.445 3.75 2.115 ;
      RECT 4.29 0.585 4.56 0.935 ;
      RECT 2.945 1.105 3.145 2.355 ;
      RECT 3.96 1.105 4.22 1.675 ;
      RECT 2.72 0.64 3.05 1.35 ;
      RECT 2.72 1.105 4.22 1.275 ;
      RECT 2.245 1.93 2.425 2.355 ;
      RECT 2.245 0.625 2.415 2.355 ;
      RECT 2.22 0.625 2.55 0.955 ;
      RECT 0.595 0.395 0.855 2.99 ;
      RECT 0.595 1.195 1.03 1.865 ;
  END
END scs130lp_dfxtp_4

MACRO scs130lp_dfxtp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dfxtp_lp 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.455 1.175 0.835 1.845 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.17 2.755 1.5 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4005 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.595 0.44 10.935 1.78 ;
        RECT 10.595 0.44 10.925 3 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 9.895 -0.085 10.145 0.9 ;
        RECT 8.545 -0.085 8.795 0.815 ;
        RECT 6.32 -0.085 6.57 0.685 ;
        RECT 2.26 -0.085 2.59 0.99 ;
        RECT 0.895 -0.085 1.225 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.04 3.415 ;
        RECT 10.065 1.96 10.395 3.415 ;
        RECT 8.535 2.105 8.865 3.415 ;
        RECT 5.36 2.075 5.69 3.415 ;
        RECT 2.54 2.03 2.87 3.415 ;
        RECT 0.76 2.025 1.09 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.39 1.755 9.72 2.935 ;
      RECT 8.535 1.755 9.72 1.925 ;
      RECT 10.085 1.085 10.415 1.755 ;
      RECT 9.545 1.585 10.415 1.755 ;
      RECT 8.535 1.425 8.845 1.925 ;
      RECT 9.545 0.355 9.715 2.935 ;
      RECT 9.255 0.355 9.715 0.725 ;
      RECT 7.12 2.075 7.45 2.935 ;
      RECT 7.12 2.075 8.355 2.245 ;
      RECT 8.185 0.355 8.355 2.245 ;
      RECT 9.055 0.905 9.365 1.575 ;
      RECT 8.185 0.995 9.365 1.165 ;
      RECT 7.675 0.355 8.355 0.685 ;
      RECT 6.51 1.685 6.84 2.935 ;
      RECT 5.245 1.725 8.005 1.895 ;
      RECT 7.835 0.865 8.005 1.895 ;
      RECT 5.245 1.155 5.44 1.895 ;
      RECT 7.115 0.865 8.005 1.035 ;
      RECT 7.115 0.605 7.445 1.035 ;
      RECT 7.345 1.215 7.655 1.545 ;
      RECT 4.525 0.455 4.715 1.485 ;
      RECT 6.51 1.215 7.655 1.385 ;
      RECT 6.51 0.865 6.68 1.385 ;
      RECT 5.97 0.865 6.68 1.035 ;
      RECT 5.97 0.455 6.14 1.035 ;
      RECT 4.525 0.455 6.14 0.625 ;
      RECT 4.175 1.685 4.505 2.875 ;
      RECT 4.175 1.685 5.065 1.855 ;
      RECT 4.895 0.805 5.065 1.855 ;
      RECT 4.175 0.375 4.345 2.875 ;
      RECT 5.62 1.215 6.33 1.545 ;
      RECT 5.62 0.805 5.79 1.545 ;
      RECT 4.895 0.805 5.79 0.975 ;
      RECT 3.71 0.375 4.345 0.685 ;
      RECT 3.285 1.725 3.615 2.73 ;
      RECT 3.285 1.725 3.995 1.895 ;
      RECT 3.825 0.865 3.995 1.895 ;
      RECT 3.2 0.865 3.995 1.035 ;
      RECT 3.2 0.375 3.53 1.035 ;
      RECT 1.29 2.025 1.845 3.065 ;
      RECT 1.675 0.265 1.845 3.065 ;
      RECT 1.675 1.68 3.105 1.85 ;
      RECT 2.935 1.215 3.105 1.85 ;
      RECT 2.935 1.215 3.645 1.545 ;
      RECT 1.675 0.265 2.015 0.725 ;
      RECT 0.105 2.025 0.56 3.065 ;
      RECT 0.105 0.265 0.275 3.065 ;
      RECT 1.165 0.825 1.495 1.495 ;
      RECT 0.105 0.825 1.495 0.995 ;
      RECT 0.105 0.265 0.435 0.995 ;
  END
END scs130lp_dfxtp_lp

MACRO scs130lp_diode_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_diode_0 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 0.255 0.87 3.075 ;
    END
  END DIODE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_diode_0

MACRO scs130lp_diode_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_diode_1 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7452 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 0.255 0.87 3.075 ;
    END
  END DIODE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_diode_1

MACRO scs130lp_dlclkp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlclkp_1 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.465 1.42 3.915 1.765 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.975 1.16 1.415 1.39 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.365 0.255 6.625 3.075 ;
    END
  END GCLK
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.865 -0.085 6.195 0.495 ;
        RECT 4.44 -0.085 4.77 0.515 ;
        RECT 2.79 -0.085 3.04 0.78 ;
        RECT 0.745 -0.085 1.075 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.635 1.835 6.195 3.415 ;
        RECT 4.695 2.905 5.025 3.415 ;
        RECT 2.715 2.615 3.045 3.415 ;
        RECT 0.605 2.24 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.265 1.495 5.465 2.495 ;
      RECT 5.265 1.495 6.195 1.665 ;
      RECT 5.945 0.665 6.195 1.665 ;
      RECT 5.345 0.665 6.195 0.835 ;
      RECT 5.345 0.44 5.675 0.835 ;
      RECT 3.585 2.565 3.915 3.075 ;
      RECT 0.975 2.905 2.445 3.075 ;
      RECT 2.275 2.275 2.445 3.075 ;
      RECT 0.095 1.9 0.425 3.075 ;
      RECT 0.975 1.9 1.145 3.075 ;
      RECT 3.225 2.565 3.915 2.745 ;
      RECT 3.225 2.565 5.095 2.735 ;
      RECT 4.925 1.005 5.095 2.735 ;
      RECT 3.225 2.275 3.395 2.745 ;
      RECT 2.275 2.275 3.395 2.445 ;
      RECT 0.095 1.9 1.145 2.07 ;
      RECT 0.095 0.255 0.365 3.075 ;
      RECT 4.925 1.005 5.675 1.325 ;
      RECT 2.45 0.95 2.835 1.265 ;
      RECT 0.095 0.82 0.58 1.095 ;
      RECT 0.095 0.82 1.415 0.99 ;
      RECT 1.245 0.255 1.415 0.99 ;
      RECT 2.45 0.255 2.62 1.265 ;
      RECT 0.095 0.255 0.575 1.095 ;
      RECT 1.245 0.255 2.62 0.425 ;
      RECT 3.565 2.225 4.755 2.395 ;
      RECT 4.585 0.685 4.755 2.395 ;
      RECT 1.655 1.91 2.095 2.24 ;
      RECT 1.925 0.965 2.095 2.24 ;
      RECT 3.565 1.935 3.825 2.395 ;
      RECT 1.655 1.935 3.825 2.105 ;
      RECT 1.925 0.965 2.28 1.295 ;
      RECT 3.21 0.685 4.755 0.855 ;
      RECT 3.21 0.445 3.5 0.855 ;
      RECT 4.085 1.025 4.415 2.055 ;
      RECT 2.265 1.505 3.295 1.765 ;
      RECT 3.045 1.025 3.295 1.765 ;
      RECT 3.045 1.025 4.415 1.25 ;
      RECT 1.315 2.485 2.07 2.735 ;
      RECT 1.315 1.56 1.485 2.735 ;
      RECT 1.315 1.56 1.755 1.74 ;
      RECT 1.585 0.595 1.755 1.74 ;
      RECT 0.535 1.56 1.755 1.73 ;
      RECT 0.535 1.345 0.795 1.73 ;
      RECT 1.585 0.595 2.06 0.795 ;
  END
END scs130lp_dlclkp_1

MACRO scs130lp_dlclkp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlclkp_2 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 1.46 3.845 1.76 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.96 1.13 1.335 1.39 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.365 0.255 6.59 3.075 ;
    END
  END GCLK
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 6.76 -0.085 7.055 1.095 ;
        RECT 5.865 -0.085 6.195 0.835 ;
        RECT 4.44 -0.085 4.77 0.345 ;
        RECT 2.7 -0.085 2.89 0.765 ;
        RECT 0.575 -0.085 0.905 0.495 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.785 1.815 7.055 3.415 ;
        RECT 5.775 2.045 6.195 3.415 ;
        RECT 4.66 2.685 4.99 3.415 ;
        RECT 2.56 2.685 2.89 3.415 ;
        RECT 0.64 2.97 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.215 1.705 5.55 2.495 ;
      RECT 5.215 1.705 6.195 1.875 ;
      RECT 5.945 1.005 6.195 1.875 ;
      RECT 5.345 1.005 6.195 1.175 ;
      RECT 5.345 0.71 5.675 1.175 ;
      RECT 3.335 2.345 3.665 3.075 ;
      RECT 1.15 2.905 2.165 3.075 ;
      RECT 1.995 2.345 2.165 3.075 ;
      RECT 1.15 2.63 1.32 3.075 ;
      RECT 0.12 2.63 1.32 2.8 ;
      RECT 0.12 1.91 0.46 2.8 ;
      RECT 1.995 2.345 5.045 2.515 ;
      RECT 4.875 1.345 5.045 2.515 ;
      RECT 0.12 0.255 0.29 2.8 ;
      RECT 4.875 1.345 5.735 1.535 ;
      RECT 2.36 0.935 2.73 1.265 ;
      RECT 0.12 0.665 0.455 1.095 ;
      RECT 2.36 0.265 2.53 1.265 ;
      RECT 0.12 0.665 1.255 0.835 ;
      RECT 1.075 0.265 1.255 0.835 ;
      RECT 0.12 0.255 0.405 1.095 ;
      RECT 1.075 0.265 2.53 0.435 ;
      RECT 3.07 1.985 4.705 2.175 ;
      RECT 4.535 0.525 4.705 2.175 ;
      RECT 1.42 1.93 3.4 2.11 ;
      RECT 1.42 1.9 2.025 2.11 ;
      RECT 1.855 1.015 2.025 2.11 ;
      RECT 1.855 1.015 2.19 1.265 ;
      RECT 3.07 0.525 4.705 0.695 ;
      RECT 3.07 0.485 3.4 0.695 ;
      RECT 4.035 0.875 4.365 1.815 ;
      RECT 2.205 1.475 3.235 1.76 ;
      RECT 3.025 0.875 3.235 1.76 ;
      RECT 3.025 0.875 4.365 1.065 ;
      RECT 1.545 2.28 1.825 2.735 ;
      RECT 1.07 2.28 1.825 2.45 ;
      RECT 1.07 1.56 1.24 2.45 ;
      RECT 0.46 1.56 1.675 1.73 ;
      RECT 1.505 0.605 1.675 1.73 ;
      RECT 0.46 1.345 0.72 1.73 ;
      RECT 1.505 0.605 1.955 0.845 ;
  END
END scs130lp_dlclkp_2

MACRO scs130lp_dlclkp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlclkp_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.474 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.4 1.365 3.85 1.76 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.855 1.17 1.315 1.39 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.195 1.815 7.535 3.075 ;
        RECT 7.355 0.255 7.535 3.075 ;
        RECT 6.485 1.075 7.535 1.245 ;
        RECT 7.345 0.255 7.535 1.245 ;
        RECT 6.295 1.815 7.535 1.985 ;
        RECT 6.485 0.255 6.675 1.245 ;
        RECT 6.295 1.815 6.525 3.075 ;
    END
  END GCLK
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.74 -0.085 8.035 1.095 ;
        RECT 6.845 -0.085 7.175 0.905 ;
        RECT 5.985 -0.085 6.315 0.895 ;
        RECT 4.675 -0.085 5.005 0.455 ;
        RECT 2.685 -0.085 2.945 0.78 ;
        RECT 0.55 -0.085 0.89 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.705 1.815 7.955 3.415 ;
        RECT 6.695 2.165 7.025 3.415 ;
        RECT 5.795 2.85 6.125 3.415 ;
        RECT 4.84 2.85 5.17 3.415 ;
        RECT 2.525 2.62 2.855 3.415 ;
        RECT 0.605 2.97 0.935 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.25 2.01 5.625 2.34 ;
      RECT 5.25 1.065 5.42 2.34 ;
      RECT 6.145 1.415 7.155 1.585 ;
      RECT 6.145 1.065 6.315 1.585 ;
      RECT 5.25 1.065 6.315 1.235 ;
      RECT 5.465 0.255 5.795 1.235 ;
      RECT 3.025 2.765 4.54 3.075 ;
      RECT 3.805 2.51 4.54 3.075 ;
      RECT 1.115 2.905 2.19 3.075 ;
      RECT 2.02 2.28 2.19 3.075 ;
      RECT 0.095 2.63 0.435 3.075 ;
      RECT 1.115 2.63 1.285 3.075 ;
      RECT 0.095 2.63 1.285 2.8 ;
      RECT 3.025 2.28 3.195 3.075 ;
      RECT 3.805 2.51 5.975 2.68 ;
      RECT 5.795 1.405 5.975 2.68 ;
      RECT 0.095 1.9 0.425 3.075 ;
      RECT 2.02 2.28 3.195 2.45 ;
      RECT 0.095 0.255 0.265 3.075 ;
      RECT 5.6 1.405 5.975 1.665 ;
      RECT 2.345 1.015 2.705 1.265 ;
      RECT 0.095 0.83 0.45 1.095 ;
      RECT 2.345 0.265 2.515 1.265 ;
      RECT 0.095 0.83 1.23 1 ;
      RECT 1.06 0.265 1.23 1 ;
      RECT 0.095 0.255 0.38 1.095 ;
      RECT 1.06 0.265 2.515 0.435 ;
      RECT 3.365 1.93 3.635 2.535 ;
      RECT 3.365 2.16 5.08 2.34 ;
      RECT 4.7 0.625 5.08 2.34 ;
      RECT 3.365 1.93 3.695 2.34 ;
      RECT 1.385 1.93 3.695 2.11 ;
      RECT 1.385 1.9 2.165 2.11 ;
      RECT 1.835 1.015 2.165 2.11 ;
      RECT 3.115 0.625 5.08 0.795 ;
      RECT 3.115 0.465 3.375 0.795 ;
      RECT 4.2 0.965 4.53 1.99 ;
      RECT 2.345 1.475 3.23 1.76 ;
      RECT 2.92 0.965 3.23 1.76 ;
      RECT 2.92 0.965 4.53 1.195 ;
      RECT 1.51 2.28 1.84 2.735 ;
      RECT 1.035 2.28 1.84 2.45 ;
      RECT 1.035 1.56 1.205 2.45 ;
      RECT 0.435 1.56 1.655 1.73 ;
      RECT 1.485 0.605 1.655 1.73 ;
      RECT 0.435 1.345 0.685 1.73 ;
      RECT 1.485 0.605 1.93 0.845 ;
  END
END scs130lp_dlclkp_4

MACRO scs130lp_dlclkp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlclkp_lp 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.02 1.455 5.635 1.785 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.605 1.27 2.15 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 0.3897 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.845 1.92 7.11 3.065 ;
        RECT 6.94 0.265 7.11 3.065 ;
        RECT 6.755 0.265 7.11 0.675 ;
    END
  END GCLK
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 5.965 -0.085 6.295 0.675 ;
        RECT 5.065 -0.085 5.395 1.275 ;
        RECT 3.045 -0.085 3.375 0.635 ;
        RECT 0.885 -0.085 1.215 0.535 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.24 2.665 6.57 3.415 ;
        RECT 5.18 2.315 5.51 3.415 ;
        RECT 3.18 2.865 3.51 3.415 ;
        RECT 0.675 2.33 1.005 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.71 2.315 6.04 3.065 ;
      RECT 5.71 2.315 6.655 2.485 ;
      RECT 6.485 0.905 6.655 2.485 ;
      RECT 6.485 0.905 6.76 1.575 ;
      RECT 5.885 0.905 6.215 1.365 ;
      RECT 5.885 0.905 6.76 1.075 ;
      RECT 3.78 2.155 4.14 2.335 ;
      RECT 3.97 1.325 4.14 2.335 ;
      RECT 4.67 1.965 6.275 2.135 ;
      RECT 5.945 1.545 6.275 2.135 ;
      RECT 4.67 0.505 4.84 2.135 ;
      RECT 2.92 1.325 3.25 1.715 ;
      RECT 2.92 1.325 4.14 1.495 ;
      RECT 3.81 0.265 3.98 1.495 ;
      RECT 3.81 0.505 4.84 0.675 ;
      RECT 3.81 0.265 4.195 0.675 ;
      RECT 4.65 2.315 4.98 3.065 ;
      RECT 1.64 2.515 4.98 2.685 ;
      RECT 4.32 2.315 4.98 2.685 ;
      RECT 1.64 1.065 1.81 2.685 ;
      RECT 4.32 0.895 4.49 2.685 ;
      RECT 1.64 1.45 2.71 1.78 ;
      RECT 1.48 1.065 1.81 1.45 ;
      RECT 0.445 1.065 1.81 1.395 ;
      RECT 4.16 0.895 4.49 1.145 ;
      RECT 2.075 2.075 3.6 2.335 ;
      RECT 3.43 1.675 3.6 2.335 ;
      RECT 3.43 1.675 3.79 1.935 ;
      RECT 2.6 0.815 3.63 1.145 ;
      RECT 2.6 0.265 2.77 1.145 ;
      RECT 1.785 0.265 2.77 0.535 ;
      RECT 0.095 2.33 0.475 3.065 ;
      RECT 0.095 0.265 0.265 3.065 ;
      RECT 2.09 0.715 2.42 1.095 ;
      RECT 0.095 0.715 2.42 0.885 ;
      RECT 0.095 0.265 0.425 0.885 ;
  END
END scs130lp_dlclkp_lp

MACRO scs130lp_dlrbn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrbn_1 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.21 2.255 1.58 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.48 2.175 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5733 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.765 1.815 9.515 3.075 ;
        RECT 9.055 0.29 9.515 3.075 ;
        RECT 9.01 0.29 9.515 1.14 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.835 1.85 8.115 3.075 ;
        RECT 7.835 0.595 8.095 3.075 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.905 1.17 6.65 1.76 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 8.605 -0.085 8.84 1.09 ;
        RECT 6.39 -0.085 6.72 0.66 ;
        RECT 4.685 -0.085 4.92 0.72 ;
        RECT 1.8 -0.085 2.02 1.04 ;
        RECT 0.105 -0.085 0.435 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 8.285 1.815 8.545 3.415 ;
        RECT 6.455 1.93 6.81 3.415 ;
        RECT 5.56 2.27 5.89 3.415 ;
        RECT 4.4 2.195 4.73 3.415 ;
        RECT 1.905 2.435 2.245 3.415 ;
        RECT 1.835 1.775 2.165 2.605 ;
        RECT 0.15 2.345 0.48 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.06 1.93 6.285 3.075 ;
      RECT 5.425 1.93 6.285 2.1 ;
      RECT 5.425 1.355 5.735 2.1 ;
      RECT 5.54 0.255 5.735 2.1 ;
      RECT 4.775 1.355 5.735 1.685 ;
      RECT 8.265 1.26 8.885 1.59 ;
      RECT 6.82 0.83 7.08 1.515 ;
      RECT 6.9 0.255 7.08 1.515 ;
      RECT 8.265 0.255 8.435 1.59 ;
      RECT 5.54 0.83 7.08 1 ;
      RECT 5.54 0.255 5.93 1 ;
      RECT 6.9 0.255 8.435 0.425 ;
      RECT 6.98 1.815 7.665 2.485 ;
      RECT 7.395 0.705 7.665 2.485 ;
      RECT 7.25 0.705 7.665 1.035 ;
      RECT 3.555 0.945 5.37 1.175 ;
      RECT 5.14 0.39 5.37 1.175 ;
      RECT 4.925 1.855 5.255 2.26 ;
      RECT 3.135 1.855 3.355 2.26 ;
      RECT 3.135 1.855 5.255 2.025 ;
      RECT 2.765 0.605 2.99 1.21 ;
      RECT 2.765 0.605 4.515 0.775 ;
      RECT 4.29 0.39 4.515 0.775 ;
      RECT 2.425 1.775 2.625 2.445 ;
      RECT 2.425 0.265 2.595 2.445 ;
      RECT 2.19 0.71 2.595 1.04 ;
      RECT 2.425 0.265 4.12 0.435 ;
      RECT 3.345 2.43 3.675 3.075 ;
      RECT 2.795 2.43 3.675 2.71 ;
      RECT 3.61 2.195 3.94 2.705 ;
      RECT 2.795 1.515 2.965 2.71 ;
      RECT 2.795 1.515 3.385 1.685 ;
      RECT 3.16 0.945 3.385 1.685 ;
      RECT 0.66 2.775 1.735 3.075 ;
      RECT 0.66 1.505 0.85 3.075 ;
      RECT 0.66 1.505 1.065 2.175 ;
      RECT 0.66 0.34 0.83 3.075 ;
      RECT 0.605 0.34 0.83 0.67 ;
      RECT 1.245 1.775 1.66 2.455 ;
      RECT 1.245 0.76 1.415 2.455 ;
      RECT 1.245 0.76 1.63 1.04 ;
      RECT 1.035 0.28 1.365 1.03 ;
  END
END scs130lp_dlrbn_1

MACRO scs130lp_dlrbn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrbn_2 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.575 1.21 2.03 1.75 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.47 2.49 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.795 0.34 7.065 1.155 ;
        RECT 6.795 1.815 7.055 2.155 ;
        RECT 6.795 0.34 6.965 2.155 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.795 0.255 9.035 3.075 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.915 1.21 6.625 2.155 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 9.205 -0.085 9.495 1.13 ;
        RECT 8.285 -0.085 8.615 0.715 ;
        RECT 7.285 -0.085 7.595 1.155 ;
        RECT 6.295 -0.085 6.625 1.04 ;
        RECT 4.545 -0.085 4.765 0.765 ;
        RECT 1.575 -0.085 1.795 1.04 ;
        RECT 0.11 -0.085 0.44 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 9.205 1.815 9.495 3.415 ;
        RECT 8.305 2.105 8.625 3.415 ;
        RECT 7.225 2.665 7.555 3.415 ;
        RECT 6.345 2.665 6.675 3.415 ;
        RECT 5.525 2.665 5.765 3.415 ;
        RECT 4.31 2.115 4.64 3.415 ;
        RECT 1.69 1.92 1.94 3.415 ;
        RECT 0.14 2.66 0.47 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 7.75 1.755 8.02 2.485 ;
      RECT 7.75 1.755 8.615 1.925 ;
      RECT 8.365 0.885 8.615 1.925 ;
      RECT 7.765 0.885 8.615 1.115 ;
      RECT 5.935 2.325 6.175 3.075 ;
      RECT 5.565 2.325 7.58 2.495 ;
      RECT 7.225 1.405 7.58 2.495 ;
      RECT 5.565 0.28 5.735 2.495 ;
      RECT 4.71 1.325 5.735 1.605 ;
      RECT 5.465 0.28 5.735 1.605 ;
      RECT 7.145 1.405 8.155 1.575 ;
      RECT 3.44 0.965 5.235 1.155 ;
      RECT 4.935 0.455 5.235 1.155 ;
      RECT 4.835 1.775 5.165 2.17 ;
      RECT 3.04 1.775 3.32 2.115 ;
      RECT 3.04 1.775 5.165 1.945 ;
      RECT 2.55 0.615 2.76 1.15 ;
      RECT 2.55 0.615 4.375 0.795 ;
      RECT 3.8 2.285 4.13 3.025 ;
      RECT 2.7 2.285 4.13 2.595 ;
      RECT 3.515 2.115 3.845 2.595 ;
      RECT 2.7 1.425 2.87 2.595 ;
      RECT 2.7 1.425 3.26 1.595 ;
      RECT 2.93 0.965 3.26 1.595 ;
      RECT 2.13 1.92 2.46 2.445 ;
      RECT 2.2 1.775 2.46 2.445 ;
      RECT 2.2 0.7 2.38 2.445 ;
      RECT 2.21 0.255 2.38 2.445 ;
      RECT 1.965 0.7 2.38 1.04 ;
      RECT 2.21 0.255 3.955 0.445 ;
      RECT 0.64 2.775 1.52 3.075 ;
      RECT 0.64 1.25 0.9 3.075 ;
      RECT 0.64 1.25 1.055 1.58 ;
      RECT 0.64 0.7 0.82 3.075 ;
      RECT 0.61 0.7 0.82 1.03 ;
      RECT 1.115 1.775 1.405 2.445 ;
      RECT 1.235 0.28 1.405 2.445 ;
      RECT 1.075 0.28 1.405 1.08 ;
      RECT 0.81 0.28 1.405 0.45 ;
  END
END scs130lp_dlrbn_2

MACRO scs130lp_dlrbn_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrbn_lp 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.09 0.835 1.78 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 0.96 1.5 1.78 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.705 1.18 8.055 3.065 ;
        RECT 7.51 0.745 7.875 1.205 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.38 1.85 9.97 2.89 ;
        RECT 9.8 0.36 9.97 2.89 ;
        RECT 9.64 0.36 9.97 0.82 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.335 1.605 6.665 2.52 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.85 -0.085 9.18 0.82 ;
        RECT 6.72 -0.085 7.05 1.075 ;
        RECT 5.345 -0.085 5.675 0.425 ;
        RECT 3.045 -0.085 3.375 0.675 ;
        RECT 0.905 -0.085 1.235 0.78 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.85 1.85 9.18 3.415 ;
        RECT 7.195 2.075 7.525 3.415 ;
        RECT 4.985 2.385 5.315 3.415 ;
        RECT 3.015 2.405 3.265 3.415 ;
        RECT 0.705 2.74 1.035 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.235 1 8.65 2.89 ;
      RECT 9.155 1 9.485 1.67 ;
      RECT 8.235 1 9.485 1.17 ;
      RECT 8.235 0.36 8.405 2.89 ;
      RECT 8.06 0.36 8.405 0.82 ;
      RECT 5.825 2.075 6.155 3.065 ;
      RECT 5.825 2.7 7.015 2.87 ;
      RECT 6.845 1.255 7.015 2.87 ;
      RECT 4.965 1.525 5.295 1.855 ;
      RECT 5.125 0.955 5.295 1.855 ;
      RECT 6.845 1.255 7.33 1.625 ;
      RECT 6.09 1.255 7.33 1.425 ;
      RECT 6.09 0.955 6.26 1.425 ;
      RECT 5.125 0.955 6.26 1.205 ;
      RECT 4.54 0.605 6.185 0.775 ;
      RECT 5.855 0.325 6.185 0.775 ;
      RECT 4.295 0.265 4.71 0.675 ;
      RECT 3.965 2.035 4.295 3.065 ;
      RECT 3.965 2.035 5.645 2.205 ;
      RECT 5.475 1.565 5.645 2.205 ;
      RECT 5.475 1.565 5.89 1.895 ;
      RECT 2.145 1.705 2.485 2.715 ;
      RECT 2.145 1.705 3.045 1.875 ;
      RECT 2.875 1.255 3.045 1.875 ;
      RECT 3.68 1.425 4.03 1.755 ;
      RECT 2.145 0.265 2.315 2.715 ;
      RECT 3.68 1.425 4.77 1.595 ;
      RECT 4.6 0.955 4.77 1.595 ;
      RECT 2.875 1.255 3.85 1.425 ;
      RECT 4.6 0.955 4.93 1.285 ;
      RECT 2.145 0.265 2.585 0.675 ;
      RECT 2.495 0.855 2.695 1.525 ;
      RECT 4.03 0.855 4.36 1.185 ;
      RECT 2.495 0.855 4.36 1.025 ;
      RECT 1.215 2.895 2.835 3.065 ;
      RECT 2.665 2.055 2.835 3.065 ;
      RECT 0.09 1.96 0.505 3 ;
      RECT 1.215 2.39 1.385 3.065 ;
      RECT 0.09 2.39 1.385 2.56 ;
      RECT 2.665 2.055 3.49 2.225 ;
      RECT 3.225 1.605 3.49 2.225 ;
      RECT 0.09 0.32 0.26 3 ;
      RECT 0.09 0.32 0.445 0.78 ;
      RECT 1.695 0.32 1.965 2.63 ;
      RECT 1.235 1.96 1.965 2.21 ;
  END
END scs130lp_dlrbn_lp

MACRO scs130lp_dlrbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrbp_1 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.45 2.345 2.12 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.995 0.885 1.755 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5649 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.62 1.74 8.075 3.075 ;
        RECT 7.815 0.26 8.075 3.075 ;
        RECT 7.605 0.26 8.075 1.06 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.75 0.26 7.055 2.155 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.945 1.21 5.47 2.12 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.225 -0.085 7.435 1.06 ;
        RECT 5.335 -0.085 5.665 0.485 ;
        RECT 4.005 -0.085 4.335 0.825 ;
        RECT 2.35 -0.085 2.645 0.94 ;
        RECT 0.715 -0.085 1.045 0.825 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.12 2.665 7.45 3.415 ;
        RECT 5.385 2.665 5.715 3.415 ;
        RECT 4.525 2.64 4.825 3.415 ;
        RECT 2.595 2.63 2.855 3.415 ;
        RECT 0.67 2.425 0.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.995 2.3 5.215 3.06 ;
      RECT 4.995 2.325 7.45 2.495 ;
      RECT 7.225 1.23 7.45 2.495 ;
      RECT 4.185 2.3 5.81 2.47 ;
      RECT 5.64 0.655 5.81 2.495 ;
      RECT 4.185 1.335 4.355 2.47 ;
      RECT 3.985 1.335 4.355 1.925 ;
      RECT 5.64 1.295 6.03 1.625 ;
      RECT 7.225 1.23 7.645 1.56 ;
      RECT 4.545 0.655 5.81 0.825 ;
      RECT 4.545 0.255 4.875 0.825 ;
      RECT 5.99 1.805 6.38 2.135 ;
      RECT 6.21 0.705 6.38 2.135 ;
      RECT 6.21 0.705 6.58 1.435 ;
      RECT 5.98 0.705 6.58 1.035 ;
      RECT 3.365 2.385 3.585 2.735 ;
      RECT 3.415 0.635 3.585 2.735 ;
      RECT 4.525 0.995 4.775 1.515 ;
      RECT 3.415 0.995 4.775 1.165 ;
      RECT 3.16 0.635 3.585 0.955 ;
      RECT 3.025 2.905 4.015 3.075 ;
      RECT 3.755 2.135 4.015 3.075 ;
      RECT 1.065 2.905 2.425 3.075 ;
      RECT 2.255 2.29 2.425 3.075 ;
      RECT 3.025 1.125 3.195 3.075 ;
      RECT 1.065 2.425 1.545 3.075 ;
      RECT 1.375 0.51 1.545 3.075 ;
      RECT 2.255 2.29 3.195 2.46 ;
      RECT 3.025 1.125 3.245 1.455 ;
      RECT 1.22 0.51 1.55 0.84 ;
      RECT 1.725 2.385 2.085 2.735 ;
      RECT 1.725 1.085 1.895 2.735 ;
      RECT 2.59 1.11 2.84 2.025 ;
      RECT 1.725 1.11 2.84 1.28 ;
      RECT 1.885 0.64 2.18 1.28 ;
      RECT 0.205 1.925 0.5 3.075 ;
      RECT 0.205 1.925 1.205 2.255 ;
      RECT 0.205 0.51 0.455 3.075 ;
      RECT 0.205 0.51 0.535 0.825 ;
  END
END scs130lp_dlrbp_1

MACRO scs130lp_dlrbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrbp_2 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.765 1.45 7.095 2.13 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.305 0.78 8.675 2.13 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.96 2.26 3.24 3.075 ;
        RECT 2.435 0.655 3.24 0.835 ;
        RECT 2.91 0.255 3.24 0.835 ;
        RECT 1.51 2.32 3.24 2.49 ;
        RECT 2.435 2.26 3.24 2.49 ;
        RECT 2.435 0.655 2.605 2.49 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5943 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 0.255 0.83 3.075 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 1.345 3.825 1.75 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 8.15 -0.085 8.415 0.61 ;
        RECT 6.57 -0.085 6.9 0.93 ;
        RECT 4.88 -0.085 5.21 0.97 ;
        RECT 3.41 -0.085 3.74 0.835 ;
        RECT 2.4 -0.085 2.73 0.465 ;
        RECT 1 -0.085 1.285 1.095 ;
        RECT 0.095 -0.085 0.385 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 8.19 2.64 8.52 3.415 ;
        RECT 6.355 2.695 6.695 3.415 ;
        RECT 4.355 2.055 4.685 3.415 ;
        RECT 3.415 2.26 3.745 3.415 ;
        RECT 2.46 2.66 2.79 3.415 ;
        RECT 1 1.815 1.29 3.415 ;
        RECT 0.095 1.815 0.385 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.69 2.3 9.025 3.065 ;
      RECT 8.845 0.28 9.025 3.065 ;
      RECT 7.955 2.3 9.025 2.47 ;
      RECT 7.955 1.585 8.135 2.47 ;
      RECT 8.585 0.28 9.025 0.61 ;
      RECT 6.865 2.81 8.02 2.98 ;
      RECT 7.615 2.64 8.02 2.98 ;
      RECT 5.115 2.785 6.165 2.955 ;
      RECT 5.995 1.125 6.165 2.955 ;
      RECT 6.865 2.355 7.035 2.98 ;
      RECT 5.115 2.055 5.445 2.955 ;
      RECT 7.615 0.28 7.785 2.98 ;
      RECT 5.995 2.355 7.035 2.525 ;
      RECT 5.965 1.125 6.165 1.455 ;
      RECT 7.615 0.28 7.98 0.61 ;
      RECT 7.205 2.3 7.435 2.64 ;
      RECT 7.265 1.1 7.435 2.64 ;
      RECT 6.335 1.1 6.595 2.025 ;
      RECT 6.335 1.1 7.435 1.27 ;
      RECT 7.07 0.64 7.33 1.27 ;
      RECT 5.625 2.275 5.825 2.615 ;
      RECT 5.625 0.64 5.795 2.615 ;
      RECT 4.25 1.185 4.545 1.535 ;
      RECT 4.25 1.185 5.795 1.355 ;
      RECT 5.625 0.64 6 0.955 ;
      RECT 3.925 1.92 4.185 3.075 ;
      RECT 3.995 1.715 4.185 3.075 ;
      RECT 3.165 1.92 4.185 2.09 ;
      RECT 3.165 1.005 3.335 2.09 ;
      RECT 3.995 1.715 5.135 1.885 ;
      RECT 4.805 1.525 5.135 1.885 ;
      RECT 2.775 1.205 3.335 1.535 ;
      RECT 3.165 1.005 4.08 1.175 ;
      RECT 4.24 0.255 4.57 1.015 ;
      RECT 3.91 0.835 4.57 1.015 ;
      RECT 1.92 0.715 2.205 2.15 ;
      RECT 1 1.3 2.205 1.63 ;
      RECT 1.875 0.715 2.205 1.63 ;
  END
END scs130lp_dlrbp_2

MACRO scs130lp_dlrbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrbp_lp 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.5 1.18 0.835 1.85 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.18 1.675 1.85 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.445 0.265 7.82 0.685 ;
        RECT 7.16 1.715 7.615 2.89 ;
        RECT 7.445 0.265 7.615 2.89 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.37 1.85 9.96 2.89 ;
        RECT 9.725 0.35 9.96 2.89 ;
        RECT 9.63 0.35 9.96 0.81 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.795 1.92 8.125 2.89 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.84 -0.085 9.17 0.81 ;
        RECT 6.7 -0.085 7.03 0.685 ;
        RECT 5.43 -0.085 5.68 0.685 ;
        RECT 3.045 -0.085 3.375 0.605 ;
        RECT 0.905 -0.085 1.235 1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.84 1.85 9.17 3.415 ;
        RECT 6.625 1.715 6.955 3.415 ;
        RECT 5.365 2.065 5.695 3.415 ;
        RECT 2.905 2.515 3.235 3.415 ;
        RECT 0.805 2.865 1.135 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.31 0.99 8.64 2.89 ;
      RECT 9.145 0.99 9.475 1.66 ;
      RECT 8.05 0.99 9.475 1.16 ;
      RECT 8.05 0.35 8.38 1.16 ;
      RECT 6.015 1.715 6.39 2.855 ;
      RECT 6.22 0.305 6.39 2.855 ;
      RECT 5.14 1.715 6.39 1.885 ;
      RECT 5.14 1.345 5.47 1.885 ;
      RECT 6.22 1.365 7.265 1.535 ;
      RECT 6.935 0.865 7.265 1.535 ;
      RECT 5.91 0.305 6.39 0.685 ;
      RECT 4.18 1.815 4.51 2.715 ;
      RECT 4.22 0.265 4.39 2.715 ;
      RECT 5.71 0.865 6.04 1.535 ;
      RECT 5.08 0.865 6.04 1.035 ;
      RECT 5.08 0.515 5.25 1.035 ;
      RECT 4.22 0.515 5.25 0.685 ;
      RECT 4.22 0.265 4.55 0.685 ;
      RECT 3.67 2.895 4.9 3.065 ;
      RECT 4.73 0.865 4.9 3.065 ;
      RECT 3.67 1.345 4 3.065 ;
      RECT 1.335 2.165 2.975 2.335 ;
      RECT 2.805 1.135 2.975 2.335 ;
      RECT 1.855 0.54 2.025 2.335 ;
      RECT 1.335 2.075 1.665 2.335 ;
      RECT 2.805 1.345 4 1.675 ;
      RECT 2.645 1.135 2.975 1.465 ;
      RECT 4.57 0.865 4.9 1.195 ;
      RECT 1.695 0.54 2.025 1 ;
      RECT 2.255 1.655 2.625 1.985 ;
      RECT 2.255 0.265 2.425 1.985 ;
      RECT 3.71 0.775 4.04 1.105 ;
      RECT 2.255 0.785 4.04 0.955 ;
      RECT 2.255 0.265 2.585 0.955 ;
      RECT 1.825 2.515 2.155 3.065 ;
      RECT 0.115 2.075 0.605 3.065 ;
      RECT 0.115 2.515 2.155 2.685 ;
      RECT 0.115 0.54 0.285 3.065 ;
      RECT 0.115 0.54 0.445 1 ;
  END
END scs130lp_dlrbp_lp

MACRO scs130lp_dlrtn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtn_1 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.375 0.815 2.005 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.8 1.325 2.005 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5733 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.075 2.64 6.635 2.97 ;
        RECT 6.37 0.255 6.635 2.97 ;
        RECT 6.09 0.255 6.635 1.095 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.425 0.84 5.74 2.13 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.59 -0.085 5.92 0.67 ;
        RECT 4.225 -0.085 4.555 0.895 ;
        RECT 2.425 -0.085 2.755 0.925 ;
        RECT 0.985 -0.085 1.205 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.575 2.64 5.905 3.415 ;
        RECT 4.295 2.285 4.915 3.415 ;
        RECT 4.65 2.025 4.915 3.415 ;
        RECT 2.5 2.655 2.83 3.415 ;
        RECT 0.685 2.515 0.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.085 2.3 5.385 3.075 ;
      RECT 5.085 2.3 6.2 2.47 ;
      RECT 5.95 1.345 6.2 2.47 ;
      RECT 5.085 0.325 5.255 3.075 ;
      RECT 4.1 1.405 4.43 2.075 ;
      RECT 4.1 1.685 5.255 1.855 ;
      RECT 5.075 0.325 5.255 1.855 ;
      RECT 4.745 0.325 5.255 0.875 ;
      RECT 3.34 2.245 3.8 2.885 ;
      RECT 3.63 0.665 3.8 2.885 ;
      RECT 4.655 1.065 4.905 1.515 ;
      RECT 3.63 1.065 4.905 1.235 ;
      RECT 3.325 0.665 3.8 0.925 ;
      RECT 1.915 0.685 2.245 2.145 ;
      RECT 3.2 1.095 3.46 2.075 ;
      RECT 1.915 1.095 3.46 1.265 ;
      RECT 2.925 0.255 3.145 1.265 ;
      RECT 2.925 0.255 3.89 0.495 ;
      RECT 1.065 2.815 2.045 2.985 ;
      RECT 1.875 2.315 2.045 2.985 ;
      RECT 0.195 2.175 0.465 2.985 ;
      RECT 1.065 2.175 1.235 2.985 ;
      RECT 1.875 2.315 2.99 2.485 ;
      RECT 2.66 1.435 2.99 2.485 ;
      RECT 0.195 2.175 1.235 2.345 ;
      RECT 0.195 0.3 0.455 2.985 ;
      RECT 1.405 2.305 1.705 2.635 ;
      RECT 1.495 0.3 1.705 2.635 ;
      RECT 1.375 0.3 1.705 0.63 ;
  END
END scs130lp_dlrtn_1

MACRO scs130lp_dlrtn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtn_2 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 0.84 0.835 1.79 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 0.84 1.295 1.79 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.905 0.255 6.115 2.145 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.26 0.685 5.52 1.515 ;
        RECT 4.945 0.685 5.52 0.855 ;
        RECT 4.945 0.375 5.185 0.855 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 6.285 -0.085 6.615 1.095 ;
        RECT 5.355 -0.085 5.685 0.515 ;
        RECT 4.005 -0.085 4.335 1 ;
        RECT 2.315 -0.085 2.645 0.955 ;
        RECT 0.7 -0.085 0.94 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 6.285 2.655 6.615 3.415 ;
        RECT 5.405 2.655 5.735 3.415 ;
        RECT 4.15 2.41 4.855 3.415 ;
        RECT 4.525 2.06 4.855 3.415 ;
        RECT 2.4 2.765 2.73 3.415 ;
        RECT 0.58 2.3 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.025 1.72 5.235 3.075 ;
      RECT 5.025 2.315 6.615 2.485 ;
      RECT 6.345 1.295 6.615 2.485 ;
      RECT 5.025 1.72 5.54 2.485 ;
      RECT 4.025 1.72 4.355 2.19 ;
      RECT 4.025 1.72 5.54 1.89 ;
      RECT 4.92 1.025 5.09 1.89 ;
      RECT 4.525 1.025 5.09 1.195 ;
      RECT 4.525 0.255 4.775 1.195 ;
      RECT 3.265 2.375 3.72 3.015 ;
      RECT 3.55 0.67 3.72 3.015 ;
      RECT 3.55 1.365 4.75 1.55 ;
      RECT 3.175 0.67 3.72 0.955 ;
      RECT 1.82 1.995 2.15 2.255 ;
      RECT 1.925 1.125 2.15 2.255 ;
      RECT 3.12 1.125 3.38 2.205 ;
      RECT 1.925 1.125 3.38 1.295 ;
      RECT 2.815 0.255 2.985 1.295 ;
      RECT 1.925 0.67 2.145 2.255 ;
      RECT 1.885 0.67 2.145 0.995 ;
      RECT 2.815 0.255 3.67 0.5 ;
      RECT 0.975 2.81 1.985 2.98 ;
      RECT 1.815 2.425 1.985 2.98 ;
      RECT 0.115 1.96 0.41 2.97 ;
      RECT 0.975 1.96 1.145 2.98 ;
      RECT 1.815 2.425 2.91 2.595 ;
      RECT 2.58 1.515 2.91 2.595 ;
      RECT 0.115 1.96 1.145 2.13 ;
      RECT 0.115 0.395 0.285 2.97 ;
      RECT 0.115 0.395 0.53 0.67 ;
      RECT 1.325 2.3 1.635 2.63 ;
      RECT 1.465 0.34 1.635 2.63 ;
      RECT 1.465 1.155 1.755 1.825 ;
      RECT 1.11 0.34 1.635 0.67 ;
  END
END scs130lp_dlrtn_2

MACRO scs130lp_dlrtn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtn_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.535 0.84 1.015 1.75 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.92 1.125 2.15 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1886 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.025 1.765 7.595 1.935 ;
        RECT 7.345 1.085 7.595 1.935 ;
        RECT 6.025 1.085 7.595 1.255 ;
        RECT 6.885 1.765 7.075 3.075 ;
        RECT 6.885 0.255 7.075 1.255 ;
        RECT 6.025 1.765 6.215 3.075 ;
        RECT 6.025 0.255 6.215 1.255 ;
        RECT 5.955 0.255 6.215 0.585 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.945 1.21 5.515 2.13 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.245 -0.085 7.575 0.915 ;
        RECT 6.385 -0.085 6.715 0.915 ;
        RECT 5.445 -0.085 5.775 0.7 ;
        RECT 4.07 -0.085 4.4 0.895 ;
        RECT 2.29 -0.085 2.62 0.875 ;
        RECT 0.795 -0.085 1.125 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.245 2.105 7.575 3.415 ;
        RECT 6.385 2.105 6.715 3.415 ;
        RECT 5.48 2.64 5.81 3.415 ;
        RECT 4.59 2.64 4.92 3.415 ;
        RECT 2.325 2.615 2.655 3.415 ;
        RECT 0.535 2.66 0.785 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.09 2.3 5.31 3.075 ;
      RECT 3.95 2.3 5.855 2.47 ;
      RECT 5.685 0.87 5.855 2.47 ;
      RECT 3.95 1.405 4.28 2.47 ;
      RECT 5.685 1.425 7.175 1.595 ;
      RECT 4.945 0.87 5.855 1.04 ;
      RECT 4.59 0.725 5.115 0.895 ;
      RECT 4.59 0.255 4.92 0.895 ;
      RECT 3.19 2.245 3.725 2.885 ;
      RECT 3.545 0.665 3.725 2.885 ;
      RECT 4.525 1.065 4.775 1.515 ;
      RECT 3.545 1.065 4.775 1.235 ;
      RECT 3.17 0.665 3.725 0.885 ;
      RECT 1.745 1.825 2.27 2.105 ;
      RECT 2.1 1.055 2.27 2.105 ;
      RECT 3.045 1.055 3.375 2.075 ;
      RECT 1.9 1.055 3.375 1.225 ;
      RECT 2.82 0.255 2.99 1.225 ;
      RECT 1.9 0.735 2.11 1.225 ;
      RECT 2.82 0.255 3.735 0.495 ;
      RECT 0.955 2.83 2.01 3 ;
      RECT 1.675 2.275 2.01 3 ;
      RECT 0.095 0.33 0.365 3 ;
      RECT 0.955 2.32 1.125 3 ;
      RECT 0.095 2.32 1.125 2.49 ;
      RECT 1.675 2.275 2.835 2.445 ;
      RECT 2.505 1.405 2.835 2.445 ;
      RECT 0.095 0.33 0.625 0.67 ;
      RECT 1.295 1.395 1.505 2.66 ;
      RECT 1.295 1.395 1.92 1.655 ;
      RECT 1.295 0.33 1.495 2.66 ;
  END
END scs130lp_dlrtn_4

MACRO scs130lp_dlrtn_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtn_lp 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.46 1.11 0.835 1.78 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 1.12 1.36 1.79 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.03 2.055 7.565 3.065 ;
        RECT 7.235 0.265 7.565 3.065 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.885 1.205 6.5 1.875 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.445 -0.085 6.775 0.675 ;
        RECT 5.175 -0.085 5.425 0.675 ;
        RECT 3.105 -0.085 3.435 0.485 ;
        RECT 0.905 -0.085 1.235 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.395 2.405 6.725 3.415 ;
        RECT 5.175 2.055 5.505 3.415 ;
        RECT 2.755 2.095 3.005 3.415 ;
        RECT 0.765 2.845 1.095 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.865 2.055 6.195 3.065 ;
      RECT 5.865 2.055 6.85 2.225 ;
      RECT 6.68 0.855 6.85 2.225 ;
      RECT 6.68 0.855 7.04 1.525 ;
      RECT 5.175 0.855 5.505 1.185 ;
      RECT 5.175 0.855 7.04 1.025 ;
      RECT 5.655 0.265 5.985 1.025 ;
      RECT 3.95 2.055 4.28 3.065 ;
      RECT 3.95 2.055 4.995 2.225 ;
      RECT 4.825 0.295 4.995 2.225 ;
      RECT 4.825 1.425 5.705 1.755 ;
      RECT 4.035 0.295 4.995 0.485 ;
      RECT 2.055 0.665 2.225 2.485 ;
      RECT 3.44 1.585 3.77 1.915 ;
      RECT 3.44 1.585 4.48 1.755 ;
      RECT 4.31 0.665 4.48 1.755 ;
      RECT 4.31 0.665 4.645 1.435 ;
      RECT 2.055 0.665 4.645 0.835 ;
      RECT 2.315 0.265 2.645 0.835 ;
      RECT 0.11 2.055 0.565 3.065 ;
      RECT 1.275 2.665 2.575 2.835 ;
      RECT 2.405 1.585 2.575 2.835 ;
      RECT 0.11 2.495 1.445 2.665 ;
      RECT 0.11 0.265 0.28 3.065 ;
      RECT 2.405 1.585 3.23 1.915 ;
      RECT 0.11 0.265 0.445 0.675 ;
      RECT 1.295 2.055 1.875 2.315 ;
      RECT 1.57 0.295 1.875 2.315 ;
      RECT 1.57 0.295 2.055 0.485 ;
      RECT 2.44 1.015 4.13 1.345 ;
  END
END scs130lp_dlrtn_lp

MACRO scs130lp_dlrtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtp_1 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.84 0.865 1.79 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 0.84 1.375 1.79 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.26 1.85 6.63 3.075 ;
        RECT 6.45 0.345 6.63 3.075 ;
        RECT 6.16 0.345 6.63 1.17 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.425 1.345 5.74 2.13 ;
        RECT 5.425 0.345 5.605 2.13 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.775 -0.085 5.99 1.17 ;
        RECT 4.345 -0.085 4.595 0.555 ;
        RECT 2.53 -0.085 2.81 0.535 ;
        RECT 0.715 -0.085 1.045 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.725 2.64 6.055 3.415 ;
        RECT 4.365 2.64 5.085 3.415 ;
        RECT 4.365 2.4 4.915 3.415 ;
        RECT 2.59 2.345 2.82 3.415 ;
        RECT 0.655 2.3 0.845 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.255 2.3 5.555 3.075 ;
      RECT 5.085 2.3 6.09 2.47 ;
      RECT 5.92 1.34 6.09 2.47 ;
      RECT 5.085 0.345 5.255 2.47 ;
      RECT 4.23 1.945 5.255 2.205 ;
      RECT 5.92 1.34 6.28 1.67 ;
      RECT 4.875 0.345 5.255 1.165 ;
      RECT 3.34 2.405 3.7 2.735 ;
      RECT 3.34 1.605 3.51 2.735 ;
      RECT 3.34 1.605 4.915 1.775 ;
      RECT 4.535 1.335 4.915 1.775 ;
      RECT 4.535 0.725 4.705 1.775 ;
      RECT 4.005 0.725 4.705 0.895 ;
      RECT 4.005 0.315 4.175 0.895 ;
      RECT 3.38 0.315 4.175 0.535 ;
      RECT 2.99 2.905 4.05 3.075 ;
      RECT 3.88 1.945 4.05 3.075 ;
      RECT 2.99 1.195 3.16 3.075 ;
      RECT 1.895 1.195 2.08 2.735 ;
      RECT 3.69 1.945 4.05 2.205 ;
      RECT 1.895 1.195 3.475 1.365 ;
      RECT 3.145 1.045 3.475 1.365 ;
      RECT 1.895 0.255 2.075 2.735 ;
      RECT 1.895 0.255 2.36 0.535 ;
      RECT 3.655 1.175 4.015 1.435 ;
      RECT 3.655 0.705 3.825 1.435 ;
      RECT 2.245 0.705 2.575 1.025 ;
      RECT 2.245 0.705 3.825 0.875 ;
      RECT 1.015 2.905 2.42 3.075 ;
      RECT 2.25 1.535 2.42 3.075 ;
      RECT 0.165 0.39 0.455 2.98 ;
      RECT 1.015 1.96 1.185 3.075 ;
      RECT 2.25 1.535 2.81 2.175 ;
      RECT 0.165 1.96 1.185 2.13 ;
      RECT 1.355 2.405 1.725 2.735 ;
      RECT 1.545 0.33 1.725 2.735 ;
      RECT 1.22 0.33 1.725 0.67 ;
  END
END scs130lp_dlrtp_1

MACRO scs130lp_dlrtp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtp_2 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.58 0.815 0.88 2.12 ;
        RECT 0.58 0.315 0.805 2.12 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.05 0.815 1.3 2.12 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6846 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.385 0.345 6.565 3.075 ;
        RECT 6.16 0.345 6.565 1.175 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.355 1.21 5.675 1.755 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 6.735 -0.085 6.985 1.225 ;
        RECT 5.605 -0.085 5.935 1.04 ;
        RECT 4.28 -0.085 4.48 0.555 ;
        RECT 2.465 -0.085 2.745 0.535 ;
        RECT 0.975 -0.085 1.175 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.735 1.815 7.075 3.415 ;
        RECT 5.75 2.265 6.08 3.415 ;
        RECT 4.29 2.63 5.05 3.415 ;
        RECT 4.29 2.44 4.785 3.415 ;
        RECT 2.645 2.395 2.835 3.415 ;
        RECT 0.6 2.695 0.85 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.22 1.925 5.47 3.075 ;
      RECT 4.955 1.925 5.47 2.46 ;
      RECT 4.24 1.905 5.125 2.235 ;
      RECT 4.24 1.925 6.215 2.095 ;
      RECT 5.965 1.345 6.215 2.095 ;
      RECT 4.955 0.345 5.125 2.46 ;
      RECT 4.81 0.345 5.125 1.165 ;
      RECT 3.355 2.405 3.72 2.655 ;
      RECT 3.355 1.555 3.525 2.655 ;
      RECT 3.355 1.555 4.775 1.725 ;
      RECT 4.47 1.335 4.775 1.725 ;
      RECT 4.47 0.725 4.64 1.725 ;
      RECT 3.94 0.725 4.64 0.895 ;
      RECT 3.94 0.255 4.11 0.895 ;
      RECT 3.315 0.255 4.11 0.535 ;
      RECT 3.005 2.825 4.07 2.995 ;
      RECT 3.9 1.905 4.07 2.995 ;
      RECT 3.005 1.045 3.175 2.995 ;
      RECT 1.885 1.535 2.135 2.715 ;
      RECT 3.705 1.905 4.07 2.235 ;
      RECT 1.82 1.535 3.175 1.705 ;
      RECT 1.82 0.255 2.01 1.705 ;
      RECT 3.005 1.045 3.41 1.305 ;
      RECT 1.82 0.255 2.295 0.535 ;
      RECT 3.59 1.125 3.95 1.385 ;
      RECT 2.18 0.705 2.51 1.365 ;
      RECT 3.59 0.705 3.76 1.385 ;
      RECT 2.18 0.705 3.76 0.875 ;
      RECT 1.02 2.885 2.475 3.055 ;
      RECT 2.305 1.895 2.475 3.055 ;
      RECT 0.16 2.355 0.43 3.025 ;
      RECT 1.02 2.355 1.19 3.055 ;
      RECT 0.16 2.355 1.19 2.525 ;
      RECT 0.16 0.315 0.41 3.025 ;
      RECT 2.305 1.895 2.835 2.225 ;
      RECT 1.36 2.355 1.715 2.715 ;
      RECT 1.48 1.885 1.715 2.715 ;
      RECT 1.48 0.33 1.65 2.715 ;
      RECT 1.425 0.33 1.65 0.66 ;
  END
END scs130lp_dlrtp_2

MACRO scs130lp_dlrtp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtp_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.84 0.875 2.13 ;
        RECT 0.625 0.47 0.805 2.13 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 0.84 1.375 2.13 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.395 1.745 8.075 1.915 ;
        RECT 7.345 1.105 8.075 1.915 ;
        RECT 6.4 1.065 7.495 1.235 ;
        RECT 7.345 1.055 7.495 1.915 ;
        RECT 7.225 0.345 7.45 1.235 ;
        RECT 7.255 1.745 7.445 3.075 ;
        RECT 6.4 0.355 6.625 1.235 ;
        RECT 6.395 1.745 6.585 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.315 1.21 5.885 2.12 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.62 -0.085 7.95 0.935 ;
        RECT 6.795 -0.085 7.055 0.895 ;
        RECT 5.9 -0.085 6.23 0.7 ;
        RECT 4.435 -0.085 4.74 0.555 ;
        RECT 2.54 -0.085 2.87 0.485 ;
        RECT 0.975 -0.085 1.165 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.615 2.085 7.945 3.415 ;
        RECT 6.755 2.085 7.085 3.415 ;
        RECT 5.85 2.63 6.18 3.415 ;
        RECT 4.96 2.63 5.29 3.415 ;
        RECT 2.835 2.335 3.035 3.415 ;
        RECT 0.645 2.64 0.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.46 2.29 5.66 3.075 ;
      RECT 4.38 2.29 6.225 2.46 ;
      RECT 6.055 0.87 6.225 2.46 ;
      RECT 4.38 1.855 4.695 2.46 ;
      RECT 6.055 1.405 7.175 1.575 ;
      RECT 6.055 0.87 6.23 1.575 ;
      RECT 5.02 0.87 6.23 1.04 ;
      RECT 5.02 0.36 5.23 1.04 ;
      RECT 3.555 2.385 3.87 2.715 ;
      RECT 3.555 1.475 3.725 2.715 ;
      RECT 3.555 1.475 5.055 1.645 ;
      RECT 4.255 1.315 5.055 1.645 ;
      RECT 4.255 0.725 4.425 1.645 ;
      RECT 4.085 0.265 4.265 0.895 ;
      RECT 3.44 0.265 4.265 0.485 ;
      RECT 3.205 2.885 4.21 3.075 ;
      RECT 4.04 1.855 4.21 3.075 ;
      RECT 3.205 0.995 3.375 3.075 ;
      RECT 2.03 2.405 2.325 2.735 ;
      RECT 2.145 1.195 2.325 2.735 ;
      RECT 3.895 1.855 4.21 2.185 ;
      RECT 1.895 1.195 3.375 1.365 ;
      RECT 3.205 0.995 3.535 1.255 ;
      RECT 1.895 0.285 2.065 1.365 ;
      RECT 1.895 0.285 2.36 0.485 ;
      RECT 3.745 1.065 4.075 1.305 ;
      RECT 3.745 0.655 3.915 1.305 ;
      RECT 2.245 0.655 2.575 1.025 ;
      RECT 2.245 0.655 3.915 0.825 ;
      RECT 1.065 2.905 2.665 3.075 ;
      RECT 2.495 1.535 2.665 3.075 ;
      RECT 0.205 2.3 0.475 2.97 ;
      RECT 1.065 2.3 1.235 3.075 ;
      RECT 0.205 2.3 1.235 2.47 ;
      RECT 0.205 0.395 0.455 2.97 ;
      RECT 2.495 1.535 3.025 2.165 ;
      RECT 1.405 2.3 1.715 2.665 ;
      RECT 1.545 0.395 1.715 2.665 ;
      RECT 1.545 1.535 1.965 2.155 ;
      RECT 1.335 0.395 1.715 0.67 ;
  END
END scs130lp_dlrtp_4

MACRO scs130lp_dlrtp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtp_lp 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.08 2.97 1.41 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 2.15 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6195 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.11 0.265 10.44 3.065 ;
        RECT 9.645 0.265 10.44 1.095 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.79 1.345 8.12 1.78 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 7.915 -0.085 8.245 0.465 ;
        RECT 5.655 -0.085 5.985 0.815 ;
        RECT 2.375 -0.085 2.705 0.715 ;
        RECT 0.115 -0.085 0.445 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.29 2.165 9.62 3.415 ;
        RECT 7.59 2.675 7.84 3.415 ;
        RECT 5.945 2.045 6.275 3.415 ;
        RECT 2.405 1.94 2.735 3.415 ;
        RECT 0.115 2.33 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.3 1.815 8.63 2.145 ;
      RECT 8.3 1.815 9.245 1.985 ;
      RECT 9.075 0.645 9.245 1.985 ;
      RECT 9.075 1.185 9.465 1.515 ;
      RECT 6.675 0.265 7.005 0.935 ;
      RECT 6.675 0.645 9.245 0.815 ;
      RECT 6.675 0.265 7.425 0.815 ;
      RECT 8.81 2.165 9.06 3.065 ;
      RECT 7.08 1.815 7.41 3.065 ;
      RECT 7.08 2.325 9.06 2.495 ;
      RECT 4.49 1.345 4.74 2.205 ;
      RECT 8.565 0.995 8.895 1.625 ;
      RECT 4.49 1.345 7.55 1.515 ;
      RECT 7.22 0.995 7.55 1.515 ;
      RECT 4.835 0.615 5.085 1.515 ;
      RECT 7.22 0.995 8.895 1.165 ;
      RECT 6.49 1.695 6.82 2.375 ;
      RECT 4.955 1.695 5.285 2.155 ;
      RECT 4.955 1.695 6.82 1.865 ;
      RECT 5.265 0.995 6.495 1.165 ;
      RECT 6.165 0.485 6.495 1.165 ;
      RECT 5.265 0.265 5.435 1.165 ;
      RECT 4.29 0.265 4.62 0.945 ;
      RECT 4.29 0.265 5.435 0.435 ;
      RECT 3.98 2.385 5.765 2.555 ;
      RECT 5.515 2.045 5.765 2.555 ;
      RECT 3.98 1.755 4.31 2.555 ;
      RECT 3.5 2.735 5.765 3.065 ;
      RECT 3.5 1.405 3.75 3.065 ;
      RECT 3.5 1.405 4.11 1.575 ;
      RECT 3.94 0.545 4.11 1.575 ;
      RECT 3.165 0.545 4.11 0.715 ;
      RECT 3.165 0.345 3.495 0.715 ;
      RECT 0.905 2.33 1.235 3.01 ;
      RECT 1.065 0.265 1.235 3.01 ;
      RECT 1.98 1.59 3.32 1.76 ;
      RECT 3.15 0.895 3.32 1.76 ;
      RECT 1.98 0.895 2.31 1.76 ;
      RECT 3.15 0.895 3.76 1.225 ;
      RECT 1.98 0.265 2.15 1.76 ;
      RECT 0.905 0.265 1.235 0.725 ;
      RECT 0.905 0.265 2.15 0.435 ;
      RECT 1.465 0.615 1.8 3.065 ;
  END
END scs130lp_dlrtp_lp

MACRO scs130lp_dlrtp_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlrtp_lp2 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.195 0.805 1.865 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.495 1.285 1.825 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.005 2.075 7.565 3.065 ;
        RECT 7.315 0.265 7.565 3.065 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.25 1.225 6.595 1.895 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.445 -0.085 6.775 0.695 ;
        RECT 5.05 -0.085 5.38 0.675 ;
        RECT 2.835 -0.085 3.165 0.545 ;
        RECT 0.935 -0.085 1.265 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.43 2.075 6.76 3.415 ;
        RECT 5.29 2.075 5.62 3.415 ;
        RECT 2.615 2.665 2.945 3.415 ;
        RECT 0.645 2.785 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.9 2.075 6.23 3.065 ;
      RECT 5.9 0.265 6.07 3.065 ;
      RECT 6.775 0.875 7.105 1.545 ;
      RECT 5.29 0.855 5.62 1.185 ;
      RECT 5.9 0.875 7.105 1.045 ;
      RECT 5.625 0.265 6.07 1.025 ;
      RECT 5.29 0.855 6.07 1.025 ;
      RECT 4.165 2.195 4.495 3.065 ;
      RECT 4.165 2.195 5.11 2.365 ;
      RECT 4.94 0.855 5.11 2.365 ;
      RECT 4.94 1.425 5.72 1.755 ;
      RECT 4.7 0.855 5.11 1.025 ;
      RECT 4.7 0.295 4.87 1.025 ;
      RECT 3.795 0.295 4.87 0.545 ;
      RECT 2.165 2.315 2.415 3.065 ;
      RECT 2.165 2.315 3.985 2.485 ;
      RECT 3.815 1.845 3.985 2.485 ;
      RECT 3.815 1.845 4.76 2.015 ;
      RECT 4.35 1.265 4.76 2.015 ;
      RECT 4.35 0.925 4.52 2.015 ;
      RECT 3.57 0.925 4.52 1.095 ;
      RECT 3.57 0.725 3.86 1.095 ;
      RECT 2.315 0.725 3.86 0.895 ;
      RECT 2.315 0.265 2.485 0.895 ;
      RECT 2.045 0.265 2.485 0.675 ;
      RECT 1.255 2.005 1.635 2.255 ;
      RECT 1.465 1.455 1.635 2.255 ;
      RECT 1.465 1.455 2.54 1.785 ;
      RECT 2.37 1.075 2.54 1.785 ;
      RECT 3.22 1.335 4.17 1.665 ;
      RECT 1.805 0.905 2.135 1.785 ;
      RECT 3.22 1.075 3.39 1.665 ;
      RECT 2.37 1.075 3.39 1.245 ;
      RECT 0.09 2.075 0.445 3.065 ;
      RECT 0.09 2.435 1.985 2.605 ;
      RECT 1.815 1.965 1.985 2.605 ;
      RECT 1.815 1.965 3.04 2.135 ;
      RECT 2.75 1.425 3.04 2.135 ;
      RECT 0.09 0.59 0.26 3.065 ;
      RECT 0.09 0.59 0.445 1.015 ;
  END
END scs130lp_dlrtp_lp2

MACRO scs130lp_dlxbn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxbn_1 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.455 1.205 0.9 1.875 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 0.255 1.775 0.675 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.805 0.255 8.065 3.075 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.59 1.805 7.125 3.075 ;
        RECT 6.785 0.995 7.125 3.075 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.305 -0.085 7.635 0.485 ;
        RECT 6.065 -0.085 6.275 0.905 ;
        RECT 4.29 -0.085 4.6 1.095 ;
        RECT 2.315 -0.085 2.645 0.505 ;
        RECT 0.675 -0.085 0.89 1.035 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.305 1.815 7.635 3.415 ;
        RECT 6.09 1.805 6.35 3.415 ;
        RECT 4.155 2.425 4.755 3.415 ;
        RECT 2.35 2.825 2.68 3.415 ;
        RECT 0.64 2.455 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.925 1.925 5.24 3.075 ;
      RECT 4.1 1.925 5.24 2.255 ;
      RECT 5.015 0.255 5.195 3.075 ;
      RECT 7.295 0.655 7.625 1.515 ;
      RECT 5.725 1.075 6.615 1.245 ;
      RECT 6.445 0.655 6.615 1.245 ;
      RECT 4.77 0.255 5.195 1.095 ;
      RECT 5.725 0.255 5.895 1.245 ;
      RECT 6.445 0.655 7.625 0.825 ;
      RECT 4.77 0.255 5.895 0.675 ;
      RECT 5.59 1.415 5.92 2.485 ;
      RECT 5.59 1.415 6.615 1.635 ;
      RECT 5.365 1.415 6.615 1.585 ;
      RECT 5.365 0.855 5.555 1.585 ;
      RECT 3.315 2.395 3.73 3.065 ;
      RECT 3.315 2.395 3.93 2.565 ;
      RECT 3.76 1.575 3.93 2.565 ;
      RECT 3.76 1.575 4.12 1.745 ;
      RECT 3.95 0.275 4.12 1.745 ;
      RECT 4.585 1.275 4.845 1.605 ;
      RECT 3.95 1.275 4.845 1.445 ;
      RECT 3.165 0.275 4.12 0.485 ;
      RECT 1.775 2.455 2.105 3.075 ;
      RECT 1.775 2.455 3.145 2.635 ;
      RECT 2.975 1.925 3.145 2.635 ;
      RECT 2.975 1.925 3.58 2.225 ;
      RECT 3.41 0.675 3.58 2.225 ;
      RECT 3.41 0.675 3.78 1.095 ;
      RECT 1.945 0.675 3.78 0.845 ;
      RECT 1.945 0.285 2.135 0.845 ;
      RECT 1.07 1.195 2.2 1.945 ;
      RECT 2.98 1.015 3.24 1.685 ;
      RECT 1.07 1.195 3.24 1.365 ;
      RECT 1.07 0.845 1.515 1.945 ;
      RECT 0.105 2.045 0.46 2.695 ;
      RECT 0.105 2.115 2.77 2.285 ;
      RECT 2.44 1.585 2.77 2.285 ;
      RECT 0.105 0.695 0.275 2.695 ;
      RECT 0.105 0.695 0.505 1.035 ;
  END
END scs130lp_dlxbn_1

MACRO scs130lp_dlxbn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxbn_2 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.45 1.21 0.91 1.88 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.32 1.61 0.65 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.705 0.655 8.045 2.135 ;
        RECT 7.775 0.33 8.045 2.135 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.765 0.965 7.095 3.075 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.64 0.085 ;
        RECT 8.215 -0.085 8.545 1.125 ;
        RECT 7.275 -0.085 7.605 0.455 ;
        RECT 6.22 -0.085 6.55 0.455 ;
        RECT 4.265 -0.085 4.595 0.885 ;
        RECT 2.22 -0.085 2.55 0.455 ;
        RECT 0.655 -0.085 0.875 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.64 3.415 ;
        RECT 8.135 2.645 8.465 3.415 ;
        RECT 7.265 2.645 7.595 3.415 ;
        RECT 6.135 1.795 6.585 3.415 ;
        RECT 4.245 2.235 4.835 3.415 ;
        RECT 2.34 2.835 2.67 3.415 ;
        RECT 0.685 2.495 1.015 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.005 1.795 5.265 3.075 ;
      RECT 5.085 0.255 5.265 3.075 ;
      RECT 7.275 2.305 8.49 2.475 ;
      RECT 8.225 1.295 8.49 2.475 ;
      RECT 7.275 0.625 7.445 2.475 ;
      RECT 4.13 1.795 5.265 2.065 ;
      RECT 4.13 1.395 4.335 2.065 ;
      RECT 4.845 0.255 5.265 1.125 ;
      RECT 5.71 0.625 7.445 0.795 ;
      RECT 5.71 0.255 6.04 0.795 ;
      RECT 4.845 0.255 6.04 0.455 ;
      RECT 5.67 0.965 5.965 2.485 ;
      RECT 5.67 1.295 6.585 1.625 ;
      RECT 5.67 0.965 6 1.625 ;
      RECT 3.28 2.39 3.61 3.075 ;
      RECT 3.28 2.39 3.96 2.56 ;
      RECT 3.79 0.255 3.96 2.56 ;
      RECT 4.505 1.295 4.915 1.625 ;
      RECT 4.505 1.055 4.675 1.625 ;
      RECT 3.79 1.055 4.675 1.225 ;
      RECT 3.15 0.255 3.96 0.455 ;
      RECT 1.77 2.495 2.1 3.075 ;
      RECT 1.77 2.495 3.1 2.665 ;
      RECT 2.93 1.965 3.1 2.665 ;
      RECT 2.93 1.965 3.62 2.22 ;
      RECT 3.38 0.625 3.62 2.22 ;
      RECT 1.78 0.625 3.62 0.795 ;
      RECT 1.78 0.28 2.05 0.795 ;
      RECT 1.23 0.965 1.56 1.985 ;
      RECT 1.23 0.965 2.185 1.955 ;
      RECT 2.935 0.965 3.21 1.755 ;
      RECT 1.23 0.965 3.21 1.375 ;
      RECT 1.045 0.82 1.4 1.09 ;
      RECT 0.11 2.06 0.515 2.73 ;
      RECT 0.11 2.155 2.76 2.325 ;
      RECT 2.435 1.625 2.76 2.325 ;
      RECT 0.11 2.06 0.53 2.325 ;
      RECT 0.11 0.7 0.28 2.73 ;
      RECT 0.11 0.7 0.485 1.04 ;
  END
END scs130lp_dlxbn_2

MACRO scs130lp_dlxbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxbp_1 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.455 0.84 0.915 1.51 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 0.255 1.775 1.115 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.35 1.815 5.665 3.075 ;
        RECT 5.495 0.255 5.665 3.075 ;
        RECT 5.35 0.255 5.665 1.095 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.325 0.375 7.595 3.075 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.825 -0.085 7.155 1.175 ;
        RECT 5.835 -0.085 6.135 1.17 ;
        RECT 4.075 -0.085 4.53 0.805 ;
        RECT 2.34 -0.085 2.67 0.575 ;
        RECT 0.66 -0.085 0.915 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.825 1.845 7.155 3.415 ;
        RECT 5.835 1.815 6.135 3.415 ;
        RECT 4.02 2.355 4.73 3.415 ;
        RECT 4.4 2.115 4.73 3.415 ;
        RECT 2.295 2.765 2.555 3.415 ;
        RECT 0.725 2.075 0.985 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.305 0.79 6.635 2.495 ;
      RECT 6.305 1.345 7.155 1.675 ;
      RECT 4.9 1.775 5.16 3.055 ;
      RECT 4.935 1.265 5.16 3.055 ;
      RECT 4.02 1.315 4.21 1.985 ;
      RECT 4.02 1.775 5.16 1.945 ;
      RECT 4.935 1.265 5.315 1.595 ;
      RECT 4.935 0.255 5.105 3.055 ;
      RECT 4.72 0.255 5.105 1.005 ;
      RECT 3.015 2.765 3.85 3.075 ;
      RECT 3.68 0.665 3.85 3.075 ;
      RECT 4.38 1.185 4.755 1.515 ;
      RECT 4.38 0.975 4.55 1.515 ;
      RECT 3.68 0.975 4.55 1.145 ;
      RECT 3.48 0.665 3.85 0.835 ;
      RECT 3.48 0.275 3.65 0.835 ;
      RECT 3.225 0.275 3.65 0.575 ;
      RECT 1.795 2.425 2.125 3.075 ;
      RECT 1.795 2.425 3.51 2.595 ;
      RECT 3.31 1.015 3.51 2.595 ;
      RECT 3.05 0.745 3.31 1.185 ;
      RECT 1.945 0.745 3.31 0.915 ;
      RECT 1.945 0.28 2.135 0.915 ;
      RECT 1.155 2.075 1.45 2.755 ;
      RECT 1.155 2.075 3.14 2.255 ;
      RECT 2.89 1.365 3.14 2.255 ;
      RECT 1.085 1.365 3.14 1.535 ;
      RECT 1.085 1.285 2.32 1.535 ;
      RECT 1.99 1.085 2.32 1.535 ;
      RECT 1.085 0.365 1.36 1.535 ;
      RECT 0.26 1.705 0.555 2.755 ;
      RECT 0.085 1.705 2.68 1.905 ;
      RECT 0.085 0.34 0.285 1.905 ;
      RECT 0.085 0.34 0.49 0.67 ;
  END
END scs130lp_dlxbp_1

MACRO scs130lp_dlxbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxbp_lp 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 1.18 0.9 2.15 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.525 1.39 2.195 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5859 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.635 1.785 8.035 1.955 ;
        RECT 7.805 0.925 8.035 1.955 ;
        RECT 6.56 0.925 8.035 1.095 ;
        RECT 6.635 1.785 6.965 3.065 ;
        RECT 6.56 0.265 6.89 1.095 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5796 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.635 0.265 9.98 3.065 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.845 -0.085 9.175 1.125 ;
        RECT 7.35 -0.085 7.68 0.745 ;
        RECT 5.21 -0.085 5.54 1.095 ;
        RECT 3.145 -0.085 3.475 0.645 ;
        RECT 0.905 -0.085 1.155 0.995 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.86 1.815 9.19 3.415 ;
        RECT 7.425 2.135 7.755 3.415 ;
        RECT 5.305 2.545 5.635 3.415 ;
        RECT 3.25 2.375 3.58 3.415 ;
        RECT 0.895 2.735 1.225 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.285 1.305 8.65 2.465 ;
      RECT 8.285 1.305 9.455 1.635 ;
      RECT 8.285 0.635 8.615 2.465 ;
      RECT 6.095 1.785 6.425 3.065 ;
      RECT 6.16 1.275 6.425 3.065 ;
      RECT 4.845 2.035 6.425 2.365 ;
      RECT 6.16 1.275 7.625 1.605 ;
      RECT 6.16 0.265 6.33 3.065 ;
      RECT 6 0.265 6.33 1.095 ;
      RECT 4.07 2.575 4.4 3.035 ;
      RECT 4.07 2.575 4.625 2.745 ;
      RECT 4.455 1.685 4.625 2.745 ;
      RECT 4.455 1.685 5.03 1.855 ;
      RECT 4.86 0.295 5.03 1.855 ;
      RECT 4.86 1.275 5.97 1.605 ;
      RECT 4.045 0.295 5.03 0.645 ;
      RECT 3.945 1.335 4.275 2.165 ;
      RECT 1.92 1.525 2.17 1.855 ;
      RECT 1.92 1.525 2.96 1.845 ;
      RECT 2.63 1.175 2.96 1.845 ;
      RECT 1.92 0.615 2.09 1.855 ;
      RECT 2.63 1.335 4.52 1.505 ;
      RECT 4.35 0.825 4.52 1.505 ;
      RECT 4.35 0.825 4.68 1.155 ;
      RECT 1.725 0.615 2.09 0.995 ;
      RECT 2.38 2.035 2.71 2.715 ;
      RECT 1.57 2.035 2.71 2.205 ;
      RECT 1.57 1.175 1.74 2.205 ;
      RECT 1.375 1.175 1.74 1.345 ;
      RECT 1.375 0.265 1.545 1.345 ;
      RECT 3.81 0.825 4.14 1.155 ;
      RECT 2.325 0.825 4.14 0.995 ;
      RECT 2.325 0.265 2.655 0.995 ;
      RECT 1.375 0.265 2.655 0.435 ;
      RECT 1.405 2.895 3.07 3.065 ;
      RECT 2.9 2.025 3.07 3.065 ;
      RECT 0.105 2.385 0.435 3.065 ;
      RECT 1.405 2.385 1.575 3.065 ;
      RECT 0.105 2.385 1.575 2.555 ;
      RECT 0.105 0.535 0.275 3.065 ;
      RECT 2.9 2.025 3.735 2.195 ;
      RECT 3.405 1.865 3.735 2.195 ;
      RECT 0.105 0.535 0.445 0.995 ;
  END
END scs130lp_dlxbp_lp

MACRO scs130lp_dlxbp_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxbp_lp2 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.505 1.11 0.835 1.78 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.175 1.895 1.845 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.1 1.18 7.555 2.89 ;
        RECT 7.1 0.265 7.27 2.89 ;
        RECT 6.705 0.265 7.27 0.595 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.635 0.44 9.965 2.89 ;
        RECT 9.375 2.025 9.705 3.065 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.845 -0.085 9.175 0.9 ;
        RECT 7.495 -0.085 7.825 0.725 ;
        RECT 5.035 -0.085 5.365 0.715 ;
        RECT 3.075 -0.085 3.405 0.635 ;
        RECT 0.905 -0.085 1.235 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.845 2.025 9.175 3.415 ;
        RECT 7.755 1.815 8.085 3.415 ;
        RECT 5.49 1.985 5.82 3.415 ;
        RECT 3.03 2.535 3.36 3.415 ;
        RECT 0.755 2.885 1.085 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.285 0.265 8.615 2.855 ;
      RECT 8.285 1.59 9.195 1.76 ;
      RECT 8.865 1.09 9.195 1.76 ;
      RECT 6.275 1.635 6.605 2.985 ;
      RECT 5.49 1.635 6.76 1.805 ;
      RECT 6.59 0.775 6.76 1.805 ;
      RECT 5.49 1.475 5.81 1.805 ;
      RECT 6.59 0.895 6.92 1.565 ;
      RECT 6.145 0.775 6.76 0.945 ;
      RECT 6.145 0.265 6.475 0.945 ;
      RECT 4.13 2.815 5.31 2.985 ;
      RECT 5.14 1.125 5.31 2.985 ;
      RECT 4.13 1.945 4.46 2.985 ;
      RECT 6.02 1.125 6.35 1.455 ;
      RECT 4.685 1.125 6.35 1.295 ;
      RECT 4.685 0.335 4.855 1.295 ;
      RECT 3.975 0.335 4.855 0.635 ;
      RECT 2.285 1.675 2.75 2.005 ;
      RECT 4.64 1.475 4.96 1.805 ;
      RECT 2.285 0.265 2.455 2.005 ;
      RECT 4.335 1.475 4.96 1.645 ;
      RECT 4.335 0.815 4.505 1.645 ;
      RECT 3.74 0.815 4.505 1.145 ;
      RECT 2.285 0.815 4.505 0.985 ;
      RECT 2.285 0.265 2.615 0.985 ;
      RECT 1.215 2.185 3.1 2.355 ;
      RECT 2.93 1.165 3.1 2.355 ;
      RECT 1.215 2.025 1.695 2.355 ;
      RECT 1.215 0.825 1.385 2.355 ;
      RECT 2.93 1.425 4.155 1.755 ;
      RECT 2.77 1.165 3.1 1.495 ;
      RECT 1.215 0.825 2.055 0.995 ;
      RECT 1.725 0.265 2.055 0.995 ;
      RECT 1.95 2.535 2.28 3.065 ;
      RECT 0.115 2.025 0.475 3.065 ;
      RECT 0.115 2.535 2.28 2.705 ;
      RECT 0.115 0.265 0.285 3.065 ;
      RECT 0.115 0.265 0.445 0.725 ;
  END
END scs130lp_dlxbp_lp2

MACRO scs130lp_dlxtn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxtn_1 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.5 1.175 1.775 1.505 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.295 2.285 0.64 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.345 0.285 6.635 3.075 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.865 -0.085 6.175 1.085 ;
        RECT 4.8 -0.085 5.11 1.085 ;
        RECT 2.825 -0.085 3.155 0.485 ;
        RECT 0.72 -0.085 0.945 1.005 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.865 1.815 6.175 3.415 ;
        RECT 4.45 2.45 5.19 3.415 ;
        RECT 4.95 2.305 5.19 3.415 ;
        RECT 2.44 2.715 2.7 3.415 ;
        RECT 0.72 2.385 0.98 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.36 1.965 5.66 3.025 ;
      RECT 5.39 1.255 5.66 3.025 ;
      RECT 4.45 1.955 4.78 2.215 ;
      RECT 4.45 1.965 5.66 2.135 ;
      RECT 5.39 1.255 6.175 1.585 ;
      RECT 5.39 0.255 5.56 3.025 ;
      RECT 5.28 0.255 5.56 1.075 ;
      RECT 3.255 2.715 4.28 3.065 ;
      RECT 4.09 1.615 4.28 3.065 ;
      RECT 4.09 1.615 5.21 1.785 ;
      RECT 4.46 1.255 5.21 1.785 ;
      RECT 4.46 0.275 4.63 1.785 ;
      RECT 3.725 0.275 4.63 0.465 ;
      RECT 4.09 0.655 4.29 1.435 ;
      RECT 2.455 0.655 4.29 0.825 ;
      RECT 2.455 0.295 2.645 0.825 ;
      RECT 1.15 2.905 2.27 3.075 ;
      RECT 2.1 2.375 2.27 3.075 ;
      RECT 1.15 2.385 1.445 3.075 ;
      RECT 2.1 2.375 3.92 2.545 ;
      RECT 3.67 0.995 3.92 2.545 ;
      RECT 1.945 0.81 2.275 1.505 ;
      RECT 3.49 0.995 3.92 1.245 ;
      RECT 1.945 0.995 3.92 1.165 ;
      RECT 1.115 0.81 2.275 1.005 ;
      RECT 1.73 2.035 1.93 2.735 ;
      RECT 1.73 2.035 3.46 2.205 ;
      RECT 3.13 1.535 3.46 2.205 ;
      RECT 0.15 1.675 0.55 3.065 ;
      RECT 0.15 1.675 2.89 1.865 ;
      RECT 2.56 1.335 2.89 1.865 ;
      RECT 0.15 0.675 0.33 3.065 ;
      RECT 0.15 0.675 0.55 1.005 ;
  END
END scs130lp_dlxtn_1

MACRO scs130lp_dlxtn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxtn_2 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.49 1.2 1.855 1.49 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 0.275 2.29 0.64 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.37 0.3 6.635 3.075 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 6.805 -0.085 7.095 1.18 ;
        RECT 5.905 -0.085 6.2 1.1 ;
        RECT 4.945 -0.085 5.17 1.09 ;
        RECT 2.89 -0.085 3.22 0.475 ;
        RECT 0.675 0.81 1.005 1.025 ;
        RECT 0.675 -0.085 0.845 1.025 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.805 1.815 7.095 3.415 ;
        RECT 5.905 1.815 6.2 3.415 ;
        RECT 4.475 2.495 5.245 3.415 ;
        RECT 5.015 1.96 5.245 3.415 ;
        RECT 2.475 2.715 2.735 3.415 ;
        RECT 0.795 2.415 1.045 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.415 1.62 5.705 2.96 ;
      RECT 5.535 0.255 5.705 2.96 ;
      RECT 4.485 1.62 4.815 2.245 ;
      RECT 4.485 1.62 5.705 1.79 ;
      RECT 5.535 1.27 6.165 1.6 ;
      RECT 5.34 0.255 5.705 1.09 ;
      RECT 3.29 2.715 4.305 3.065 ;
      RECT 4.135 1.27 4.305 3.065 ;
      RECT 4.135 1.27 5.355 1.45 ;
      RECT 4.605 1.26 5.355 1.45 ;
      RECT 4.605 0.255 4.775 1.45 ;
      RECT 3.79 0.255 4.775 0.475 ;
      RECT 4.095 0.645 4.425 1.1 ;
      RECT 2.46 0.645 4.425 0.815 ;
      RECT 2.46 0.275 2.72 0.815 ;
      RECT 1.215 2.905 2.305 3.075 ;
      RECT 2.135 2.375 2.305 3.075 ;
      RECT 1.215 2.395 1.515 3.075 ;
      RECT 2.135 2.375 3.965 2.545 ;
      RECT 3.705 1.915 3.965 2.545 ;
      RECT 3.705 0.995 3.925 2.545 ;
      RECT 2.025 0.995 2.34 1.49 ;
      RECT 2.025 0.995 3.925 1.165 ;
      RECT 1.185 0.81 2.29 1.03 ;
      RECT 1.705 2.035 1.955 2.735 ;
      RECT 1.705 2.035 3.495 2.205 ;
      RECT 3.165 1.535 3.495 2.205 ;
      RECT 0.14 1.66 0.625 3.055 ;
      RECT 0.14 1.66 2.925 1.855 ;
      RECT 2.595 1.345 2.925 1.855 ;
      RECT 0.14 0.695 0.31 3.055 ;
      RECT 0.14 0.695 0.495 1.025 ;
  END
END scs130lp_dlxtn_2

MACRO scs130lp_dlxtn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxtn_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.43 1.19 1.285 1.52 ;
    END
  END D
  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 0.28 1.845 0.65 ;
    END
  END GATEN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.86 1.685 7.095 3.075 ;
        RECT 6.875 0.255 7.095 3.075 ;
        RECT 6.865 1.005 7.095 3.075 ;
        RECT 5.97 1.005 7.095 1.175 ;
        RECT 6 1.685 7.095 1.855 ;
        RECT 6 1.685 6.225 3.075 ;
        RECT 5.97 0.255 6.195 1.175 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.265 -0.085 7.495 1.095 ;
        RECT 6.365 -0.085 6.695 0.835 ;
        RECT 5.555 -0.085 5.8 1.095 ;
        RECT 4.47 -0.085 4.72 0.885 ;
        RECT 2.415 -0.085 2.745 0.455 ;
        RECT 0.64 -0.085 0.885 1.02 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.265 1.815 7.585 3.415 ;
        RECT 6.395 2.025 6.69 3.415 ;
        RECT 5.545 1.815 5.83 3.415 ;
        RECT 4.205 2.435 4.915 3.415 ;
        RECT 4.585 2.015 4.915 3.415 ;
        RECT 2.3 2.74 2.56 3.415 ;
        RECT 0.58 2.395 0.835 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.085 1.675 5.375 3.035 ;
      RECT 5.205 0.255 5.375 3.035 ;
      RECT 4.205 1.675 4.415 2.265 ;
      RECT 4.205 1.675 5.375 1.845 ;
      RECT 4.205 1.595 4.385 2.265 ;
      RECT 5.205 1.345 6.695 1.515 ;
      RECT 5.205 0.255 5.385 1.515 ;
      RECT 4.89 0.255 5.385 1.075 ;
      RECT 3.02 2.74 4.035 3.02 ;
      RECT 3.865 1.245 4.035 3.02 ;
      RECT 4.705 1.245 5.035 1.505 ;
      RECT 3.865 1.245 5.035 1.415 ;
      RECT 4.13 0.255 4.3 1.415 ;
      RECT 3.25 0.255 4.3 0.455 ;
      RECT 3.62 0.625 3.95 1.065 ;
      RECT 2.035 0.625 3.95 0.795 ;
      RECT 2.035 0.255 2.235 0.795 ;
      RECT 1.005 2.905 2.13 3.075 ;
      RECT 1.96 2.4 2.13 3.075 ;
      RECT 1.005 2.395 1.305 3.075 ;
      RECT 1.96 2.4 3.695 2.57 ;
      RECT 3.435 1.325 3.695 2.57 ;
      RECT 1.695 0.965 2.14 1.53 ;
      RECT 3.08 1.325 3.695 1.495 ;
      RECT 3.08 0.965 3.41 1.495 ;
      RECT 1.695 0.965 3.41 1.145 ;
      RECT 1.055 0.82 1.865 1.01 ;
      RECT 1.53 2.05 1.78 2.735 ;
      RECT 1.53 2.05 3.225 2.22 ;
      RECT 2.895 1.675 3.225 2.22 ;
      RECT 0.09 1.7 0.41 3.055 ;
      RECT 0.09 1.7 2.685 1.88 ;
      RECT 2.355 1.315 2.685 1.88 ;
      RECT 0.09 0.68 0.26 3.055 ;
      RECT 0.09 0.68 0.47 1.01 ;
  END
END scs130lp_dlxtn_4

MACRO scs130lp_dlxtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxtp_1 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.47 0.775 0.815 1.445 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.05 0.775 1.285 1.105 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.385 0.295 5.675 3.075 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.975 -0.085 5.215 1.095 ;
        RECT 3.9 -0.085 4.23 0.625 ;
        RECT 2.195 0.605 2.57 0.845 ;
        RECT 2.4 -0.085 2.57 0.845 ;
        RECT 0.705 -0.085 0.95 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.905 2.035 5.215 3.415 ;
        RECT 4.975 1.815 5.215 3.415 ;
        RECT 3.955 2.035 4.285 3.415 ;
        RECT 2.07 2.645 2.4 3.415 ;
        RECT 0.585 2.135 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.455 1.695 4.715 2.95 ;
      RECT 3.665 1.695 4.805 1.865 ;
      RECT 4.635 0.285 4.805 1.865 ;
      RECT 3.665 1.185 3.995 1.865 ;
      RECT 4.635 1.265 5.215 1.595 ;
      RECT 4.4 0.285 4.805 0.625 ;
      RECT 3.015 2.075 3.46 2.745 ;
      RECT 3.29 0.795 3.46 2.745 ;
      RECT 4.205 0.795 4.465 1.515 ;
      RECT 3 0.795 4.465 1.005 ;
      RECT 1.545 2.305 1.875 2.965 ;
      RECT 1.545 2.305 2.82 2.475 ;
      RECT 2.65 1.015 2.82 2.475 ;
      RECT 2.65 1.395 3.12 1.725 ;
      RECT 1.765 1.015 2.82 1.185 ;
      RECT 1.765 0.675 2.025 1.185 ;
      RECT 0.085 1.625 0.365 2.775 ;
      RECT 0.085 1.625 1.155 1.795 ;
      RECT 0.985 1.365 1.155 1.795 ;
      RECT 2.22 1.365 2.48 1.745 ;
      RECT 0.085 0.265 0.3 2.775 ;
      RECT 0.985 1.365 2.48 1.535 ;
      RECT 0.085 0.265 0.535 0.605 ;
      RECT 1.12 0.255 1.425 0.605 ;
      RECT 1.12 0.255 2.22 0.435 ;
      RECT 1.015 1.965 1.335 2.775 ;
      RECT 1.335 1.705 1.69 2.135 ;
  END
END scs130lp_dlxtp_1

MACRO scs130lp_dlxtp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxtp_lp 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.82 1.6 2.15 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 1.48 0.905 2.15 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.705 0.265 8.035 3.065 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 6.915 -0.085 7.245 1.125 ;
        RECT 5.28 -0.085 5.61 0.675 ;
        RECT 3.285 -0.085 3.615 0.545 ;
        RECT 0.905 -0.085 1.235 0.95 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 6.915 1.815 7.245 3.415 ;
        RECT 5.565 1.815 5.895 3.415 ;
        RECT 3.195 2.825 3.525 3.415 ;
        RECT 0.935 2.33 1.265 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.355 0.265 6.685 3.065 ;
      RECT 6.355 1.305 7.525 1.635 ;
      RECT 5.15 0.925 5.48 1.255 ;
      RECT 5.15 0.925 6.685 1.095 ;
      RECT 4.095 2.825 5.245 3.035 ;
      RECT 5.075 1.435 5.245 3.035 ;
      RECT 4.8 1.435 6.17 1.605 ;
      RECT 5.84 1.275 6.17 1.605 ;
      RECT 4.8 0.505 4.97 1.605 ;
      RECT 4.455 0.505 4.97 0.675 ;
      RECT 4.455 0.265 4.785 0.675 ;
      RECT 2.295 2.435 2.625 3.065 ;
      RECT 2.295 2.475 4.895 2.645 ;
      RECT 4.45 2.185 4.895 2.645 ;
      RECT 4.45 0.855 4.62 2.645 ;
      RECT 4.105 0.855 4.62 1.185 ;
      RECT 2.465 0.725 4.275 0.895 ;
      RECT 2.465 0.265 2.795 0.895 ;
      RECT 0.115 0.49 0.365 3.01 ;
      RECT 3.94 1.585 4.27 1.975 ;
      RECT 2.98 1.585 4.27 1.755 ;
      RECT 1.375 1.425 3.31 1.595 ;
      RECT 1.375 1.13 1.545 1.595 ;
      RECT 0.115 1.13 1.545 1.3 ;
      RECT 0.115 0.49 0.445 1.3 ;
      RECT 3.55 1.075 3.88 1.405 ;
      RECT 1.725 1.075 3.88 1.245 ;
      RECT 1.725 0.49 2.055 1.245 ;
      RECT 1.725 2.33 2.055 3.01 ;
      RECT 1.885 1.965 2.055 3.01 ;
      RECT 3.4 1.965 3.73 2.295 ;
      RECT 1.885 1.965 3.73 2.135 ;
  END
END scs130lp_dlxtp_lp

MACRO scs130lp_dlxtp_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlxtp_lp2 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 0.905 0.835 1.78 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.05 1.175 1.38 1.845 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.46 0.44 8.05 2.925 ;
        RECT 7.72 0.395 8.05 2.925 ;
    END
  END Q
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 6.93 -0.085 7.26 0.855 ;
        RECT 5.41 -0.085 5.74 0.675 ;
        RECT 3.045 -0.085 3.375 0.675 ;
        RECT 0.905 -0.085 1.235 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 6.93 1.885 7.26 3.415 ;
        RECT 5.41 2.075 5.74 3.415 ;
        RECT 2.85 2.935 3.18 3.415 ;
        RECT 0.645 2.805 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.14 2.075 6.565 3.065 ;
      RECT 6.395 0.265 6.565 3.065 ;
      RECT 5.41 1.705 6.565 1.875 ;
      RECT 6.395 1.035 6.965 1.705 ;
      RECT 5.41 1.205 5.675 1.875 ;
      RECT 6.395 0.265 6.7 1.705 ;
      RECT 6.37 0.265 6.7 0.675 ;
      RECT 4.305 2.075 4.635 3.065 ;
      RECT 4.305 2.075 5.23 2.245 ;
      RECT 5.06 0.295 5.23 2.245 ;
      RECT 5.885 0.855 6.215 1.525 ;
      RECT 5.06 0.855 6.215 1.025 ;
      RECT 3.945 0.295 5.23 0.585 ;
      RECT 2.24 0.265 2.57 2.405 ;
      RECT 4.61 0.765 4.88 1.895 ;
      RECT 2.24 0.915 4.88 1.085 ;
      RECT 3.71 0.765 4.88 1.085 ;
      RECT 2.24 0.265 2.585 1.085 ;
      RECT 2.75 1.265 3.08 1.935 ;
      RECT 4.07 1.265 4.4 1.665 ;
      RECT 2.75 1.265 4.4 1.435 ;
      RECT 0.115 2.025 0.445 3.065 ;
      RECT 1.155 2.585 3.65 2.755 ;
      RECT 3.32 1.615 3.65 2.755 ;
      RECT 0.115 2.455 1.325 2.625 ;
      RECT 0.115 0.265 0.285 3.065 ;
      RECT 0.115 0.265 0.445 0.725 ;
      RECT 1.175 2.025 2.025 2.275 ;
      RECT 1.695 0.265 2.025 2.275 ;
  END
END scs130lp_dlxtp_lp2

MACRO scs130lp_dlybuf4s15kapwr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s15kapwr_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 3.77 2.945 ;
      LAYER li ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s15kapwr_1

MACRO scs130lp_dlybuf4s15kapwr_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s15kapwr_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.685 4.25 2.94 ;
      LAYER li ;
        RECT 3.875 1.815 4.125 3.075 ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s15kapwr_2

MACRO scs130lp_dlybuf4s18kapwr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s18kapwr_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 3.77 2.945 ;
      LAYER li ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s18kapwr_1

MACRO scs130lp_dlybuf4s18kapwr_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s18kapwr_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 4.25 2.945 ;
      LAYER li ;
        RECT 3.875 1.815 4.125 3.075 ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s18kapwr_2

MACRO scs130lp_dlybuf4s25kapwr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s25kapwr_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 3.77 2.945 ;
      LAYER li ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s25kapwr_1

MACRO scs130lp_dlybuf4s25kapwr_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s25kapwr_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 4.25 2.945 ;
      LAYER li ;
        RECT 3.875 1.815 4.125 3.075 ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s25kapwr_2

MACRO scs130lp_dlybuf4s50kapwr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s50kapwr_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.75 3.075 ;
        RECT 3.515 0.31 3.75 3.075 ;
        RECT 3.21 0.31 3.75 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 3.77 2.945 ;
      LAYER li ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s50kapwr_1

MACRO scs130lp_dlybuf4s50kapwr_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlybuf4s50kapwr_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.55 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4704 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.23 1.815 3.705 3.075 ;
        RECT 3.515 0.31 3.705 3.075 ;
        RECT 3.21 0.31 3.705 0.64 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 4.25 2.945 ;
      LAYER li ;
        RECT 3.875 1.815 4.125 3.075 ;
        RECT 2.71 2.165 3.04 3.075 ;
        RECT 0.595 2.38 0.925 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.875 -0.085 4.125 0.645 ;
        RECT 2.71 -0.085 3.04 0.67 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.01 2.08 2.26 3.075 ;
      RECT 2.01 2.08 2.54 2.25 ;
      RECT 2.37 1.825 2.54 2.25 ;
      RECT 2.37 1.825 3.025 1.995 ;
      RECT 2.855 0.98 3.025 1.995 ;
      RECT 2.855 1.295 3.345 1.625 ;
      RECT 2.01 0.98 3.025 1.215 ;
      RECT 2.01 0.27 2.26 1.215 ;
      RECT 1.385 2.395 1.84 3.075 ;
      RECT 1.67 0.27 1.84 3.075 ;
      RECT 1.445 2.1 1.84 3.075 ;
      RECT 1.67 1.385 2.685 1.655 ;
      RECT 1.435 0.27 1.84 1.28 ;
      RECT 0.095 2.03 0.425 3.075 ;
      RECT 0.095 2.03 1.265 2.205 ;
      RECT 0.91 0.82 1.265 2.205 ;
      RECT 0.91 1.6 1.5 1.93 ;
      RECT 0.095 0.82 1.265 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlybuf4s50kapwr_2

MACRO scs130lp_dlygate4s15_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlygate4s15_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.325 1.815 3.74 3.075 ;
        RECT 3.45 0.255 3.74 3.075 ;
        RECT 3.325 0.255 3.74 1.12 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.825 -0.085 3.155 0.875 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.825 2.165 3.155 3.415 ;
        RECT 0.57 2.38 0.9 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.985 1.825 2.345 2.19 ;
      RECT 1.985 1.825 3.155 1.995 ;
      RECT 2.91 1.045 3.155 1.995 ;
      RECT 2.91 1.295 3.28 1.625 ;
      RECT 1.985 1.045 3.155 1.215 ;
      RECT 1.985 0.71 2.345 1.215 ;
      RECT 1.415 2.395 1.72 2.725 ;
      RECT 1.475 0.305 1.72 2.725 ;
      RECT 1.475 1.385 2.74 1.655 ;
      RECT 1.415 0.305 1.72 0.635 ;
      RECT 0.095 2.03 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 0.82 1.305 2.205 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlygate4s15_1

MACRO scs130lp_dlygate4s18_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlygate4s18_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.325 1.815 3.74 3.075 ;
        RECT 3.45 0.255 3.74 3.075 ;
        RECT 3.325 0.255 3.74 1.12 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.825 -0.085 3.155 0.875 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.825 2.165 3.155 3.415 ;
        RECT 0.57 2.38 0.9 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.985 1.825 2.345 2.19 ;
      RECT 1.985 1.825 3.155 1.995 ;
      RECT 2.91 1.045 3.155 1.995 ;
      RECT 2.91 1.295 3.28 1.625 ;
      RECT 1.985 1.045 3.155 1.215 ;
      RECT 1.985 0.71 2.345 1.215 ;
      RECT 1.415 2.395 1.72 2.725 ;
      RECT 1.475 0.305 1.72 2.725 ;
      RECT 1.475 1.385 2.74 1.655 ;
      RECT 1.415 0.305 1.72 0.635 ;
      RECT 0.095 2.03 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 0.82 1.305 2.205 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlygate4s18_1

MACRO scs130lp_dlygate4s50_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlygate4s50_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.325 1.815 3.74 3.075 ;
        RECT 3.45 0.255 3.74 3.075 ;
        RECT 3.325 0.255 3.74 1.12 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.825 -0.085 3.155 0.875 ;
        RECT 0.58 -0.085 0.91 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.825 2.165 3.155 3.415 ;
        RECT 0.57 2.38 0.9 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.985 1.825 2.345 2.19 ;
      RECT 1.985 1.825 3.155 1.995 ;
      RECT 2.91 1.045 3.155 1.995 ;
      RECT 2.91 1.295 3.28 1.625 ;
      RECT 1.985 1.045 3.155 1.215 ;
      RECT 1.985 0.71 2.345 1.215 ;
      RECT 1.415 2.395 1.72 2.725 ;
      RECT 1.475 0.305 1.72 2.725 ;
      RECT 1.475 1.385 2.74 1.655 ;
      RECT 1.415 0.305 1.72 0.635 ;
      RECT 0.095 2.03 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 0.82 1.305 2.205 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 1.02 ;
  END
END scs130lp_dlygate4s50_1

MACRO scs130lp_dlymetal6s2s_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlymetal6s2s_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.315 0.55 1.765 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    ANTENNADIFFAREA 0.5565 LAYER met1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.126 LAYER met1 ;
      ANTENNAMAXAREACAR 7.076984 LAYER li ;
      ANTENNAMAXAREACAR 7.076984 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 6.103175 LAYER li ;
      ANTENNAMAXSIDEAREACAR 6.103175 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 0.96 2.32 4.205 2.49 ;
        RECT 0.96 1.92 1.325 2.49 ;
      LAYER li ;
        RECT 1.18 1.315 1.99 1.605 ;
        RECT 1.06 1.835 1.35 3.075 ;
        RECT 1.18 0.255 1.35 3.075 ;
        RECT 1.085 0.255 1.35 1.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.465 -0.085 3.795 0.805 ;
        RECT 2.025 -0.085 2.355 0.805 ;
        RECT 0.585 -0.085 0.915 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.465 2.33 3.76 3.415 ;
        RECT 2.025 2.33 2.32 3.415 ;
        RECT 0.585 2.33 0.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 3.84 1.92 4.205 2.15 ;
      RECT 2.4 1.92 2.765 2.15 ;
    LAYER li ;
      RECT 3.94 1.835 4.235 3.075 ;
      RECT 4.06 0.255 4.235 3.075 ;
      RECT 3.965 0.255 4.235 1.075 ;
      RECT 2.975 1.895 3.305 2.225 ;
      RECT 2.975 1.895 3.77 2.16 ;
      RECT 3.6 0.975 3.77 2.16 ;
      RECT 3.6 1.275 3.89 1.605 ;
      RECT 2.975 0.975 3.77 1.145 ;
      RECT 2.975 0.7 3.27 1.145 ;
      RECT 2.5 1.835 2.79 3.075 ;
      RECT 2.62 0.255 2.79 3.075 ;
      RECT 2.62 1.315 3.43 1.605 ;
      RECT 2.525 0.255 2.79 1.075 ;
      RECT 1.535 1.895 1.865 2.225 ;
      RECT 1.535 1.895 2.33 2.16 ;
      RECT 2.16 0.975 2.33 2.16 ;
      RECT 2.16 1.275 2.45 1.605 ;
      RECT 1.535 0.975 2.33 1.145 ;
      RECT 1.535 0.7 1.83 1.145 ;
      RECT 0.095 1.935 0.425 2.225 ;
      RECT 0.095 1.935 0.89 2.16 ;
      RECT 0.72 0.975 0.89 2.16 ;
      RECT 0.72 1.275 1.01 1.605 ;
      RECT 0.095 0.975 0.89 1.145 ;
      RECT 0.095 0.7 0.39 1.145 ;
  END
END scs130lp_dlymetal6s2s_1

MACRO scs130lp_dlymetal6s4s_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlymetal6s4s_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.315 0.55 1.765 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    ANTENNADIFFAREA 0.5565 LAYER met1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.126 LAYER met1 ;
      ANTENNAMAXAREACAR 7.076984 LAYER li ;
      ANTENNAMAXAREACAR 7.076984 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 6.103175 LAYER li ;
      ANTENNAMAXSIDEAREACAR 6.103175 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 0.96 2.32 4.205 2.49 ;
        RECT 2.4 1.92 2.765 2.49 ;
      LAYER li ;
        RECT 2.62 1.315 3.43 1.605 ;
        RECT 2.5 1.835 2.79 3.075 ;
        RECT 2.62 0.255 2.79 3.075 ;
        RECT 2.525 0.255 2.79 1.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.465 -0.085 3.795 0.805 ;
        RECT 2.025 -0.085 2.355 0.805 ;
        RECT 0.585 -0.085 0.915 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.465 2.33 3.76 3.415 ;
        RECT 2.025 2.33 2.32 3.415 ;
        RECT 0.585 2.33 0.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 3.84 1.92 4.205 2.15 ;
      RECT 0.96 1.92 1.325 2.15 ;
    LAYER li ;
      RECT 3.94 1.835 4.235 3.075 ;
      RECT 4.06 0.255 4.235 3.075 ;
      RECT 3.965 0.255 4.235 1.075 ;
      RECT 2.975 1.895 3.305 2.225 ;
      RECT 2.975 1.895 3.77 2.16 ;
      RECT 3.6 0.975 3.77 2.16 ;
      RECT 3.6 1.275 3.89 1.605 ;
      RECT 2.975 0.975 3.77 1.145 ;
      RECT 2.975 0.7 3.27 1.145 ;
      RECT 1.535 1.895 1.865 2.225 ;
      RECT 1.535 1.895 2.33 2.16 ;
      RECT 2.16 0.975 2.33 2.16 ;
      RECT 2.16 1.275 2.45 1.605 ;
      RECT 1.535 0.975 2.33 1.145 ;
      RECT 1.535 0.7 1.83 1.145 ;
      RECT 1.06 1.835 1.35 3.075 ;
      RECT 1.18 0.255 1.35 3.075 ;
      RECT 1.18 1.315 1.99 1.605 ;
      RECT 1.085 0.255 1.35 1.075 ;
      RECT 0.095 1.935 0.425 2.225 ;
      RECT 0.095 1.935 0.89 2.16 ;
      RECT 0.72 0.975 0.89 2.16 ;
      RECT 0.72 1.275 1.01 1.605 ;
      RECT 0.095 0.975 0.89 1.145 ;
      RECT 0.095 0.7 0.39 1.145 ;
  END
END scs130lp_dlymetal6s4s_1

MACRO scs130lp_dlymetal6s6s_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_dlymetal6s6s_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.315 0.55 1.765 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    ANTENNADIFFAREA 0.5565 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.96 2.32 4.205 2.49 ;
        RECT 3.84 1.92 4.205 2.49 ;
      LAYER li ;
        RECT 3.94 1.835 4.235 3.075 ;
        RECT 4.06 0.255 4.235 3.075 ;
        RECT 3.965 0.255 4.235 1.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.465 -0.085 3.795 0.805 ;
        RECT 2.025 -0.085 2.355 0.805 ;
        RECT 0.585 -0.085 0.915 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.465 2.33 3.76 3.415 ;
        RECT 2.025 2.33 2.32 3.415 ;
        RECT 0.585 2.33 0.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 2.4 1.92 2.765 2.15 ;
      RECT 0.96 1.92 1.325 2.15 ;
    LAYER li ;
      RECT 2.975 1.895 3.305 2.225 ;
      RECT 2.975 1.895 3.77 2.16 ;
      RECT 3.6 0.975 3.77 2.16 ;
      RECT 3.6 1.275 3.89 1.605 ;
      RECT 2.975 0.975 3.77 1.145 ;
      RECT 2.975 0.7 3.27 1.145 ;
      RECT 2.5 1.835 2.79 3.075 ;
      RECT 2.62 0.255 2.79 3.075 ;
      RECT 2.62 1.315 3.43 1.605 ;
      RECT 2.525 0.255 2.79 1.075 ;
      RECT 1.535 1.895 1.865 2.225 ;
      RECT 1.535 1.895 2.33 2.16 ;
      RECT 2.16 0.975 2.33 2.16 ;
      RECT 2.16 1.275 2.45 1.605 ;
      RECT 1.535 0.975 2.33 1.145 ;
      RECT 1.535 0.7 1.83 1.145 ;
      RECT 1.06 1.835 1.35 3.075 ;
      RECT 1.18 0.255 1.35 3.075 ;
      RECT 1.18 1.315 1.99 1.605 ;
      RECT 1.085 0.255 1.35 1.075 ;
      RECT 0.095 1.935 0.425 2.225 ;
      RECT 0.095 1.935 0.89 2.16 ;
      RECT 0.72 0.975 0.89 2.16 ;
      RECT 0.72 1.275 1.01 1.605 ;
      RECT 0.095 0.975 0.89 1.145 ;
      RECT 0.095 0.7 0.39 1.145 ;
  END
END scs130lp_dlymetal6s6s_1

MACRO scs130lp_ebufn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ebufn_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.27 3.415 1.94 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.348 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.45 1.27 2.78 1.94 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.345 0.73 1.145 ;
        RECT 0.125 1.815 0.7 3.075 ;
        RECT 0.125 0.345 0.355 3.075 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.74 -0.085 3.07 1.1 ;
        RECT 1.22 -0.085 1.55 1.225 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.79 2.45 3.12 3.415 ;
        RECT 1.19 1.795 1.52 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.69 2.905 2.62 3.075 ;
      RECT 2.45 2.11 2.62 3.075 ;
      RECT 1.69 1.455 1.86 3.075 ;
      RECT 3.29 2.11 3.755 2.79 ;
      RECT 3.585 0.93 3.755 2.79 ;
      RECT 2.45 2.11 3.755 2.28 ;
      RECT 0.525 1.315 0.855 1.645 ;
      RECT 0.525 1.455 1.86 1.625 ;
      RECT 3.24 0.93 3.755 1.1 ;
      RECT 3.24 0.64 3.57 1.1 ;
      RECT 2.03 0.64 2.28 2.735 ;
      RECT 2.03 0.64 2.57 1.1 ;
      RECT 2.03 0.255 2.2 2.735 ;
      RECT 1.82 0.255 2.2 0.585 ;
  END
END scs130lp_ebufn_1

MACRO scs130lp_ebufn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ebufn_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 1.305 3.895 2.15 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.537 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.995 1.305 3.325 2.15 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5964 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.955 0.945 1.125 ;
        RECT 0.615 0.595 0.945 1.125 ;
        RECT 0.685 1.795 0.855 2.735 ;
        RECT 0.125 1.795 0.855 1.965 ;
        RECT 0.125 0.955 0.355 1.965 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.37 -0.085 3.7 1.135 ;
        RECT 1.625 -0.085 1.875 0.785 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.335 2.785 3.665 3.415 ;
        RECT 1.545 2.155 1.715 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.835 2.435 4.235 3.075 ;
      RECT 4.065 0.675 4.235 3.075 ;
      RECT 2.315 2.615 3.165 2.785 ;
      RECT 2.995 2.445 4.235 2.615 ;
      RECT 2.315 1.295 2.485 2.785 ;
      RECT 0.74 1.295 2.485 1.625 ;
      RECT 3.87 0.675 4.235 1.135 ;
      RECT 2.655 0.255 2.825 2.445 ;
      RECT 2.655 0.255 3.2 1.135 ;
      RECT 2.605 0.255 3.2 0.585 ;
      RECT 1.115 0.955 2.375 1.125 ;
      RECT 2.045 0.255 2.375 1.125 ;
      RECT 1.115 0.255 1.445 1.125 ;
      RECT 0.115 0.255 0.445 0.785 ;
      RECT 0.115 0.255 1.445 0.425 ;
      RECT 1.895 1.815 2.145 3.075 ;
      RECT 0.175 2.905 1.365 3.075 ;
      RECT 1.035 1.815 1.365 3.075 ;
      RECT 0.175 2.135 0.505 3.075 ;
      RECT 1.035 1.815 2.145 1.985 ;
  END
END scs130lp_ebufn_2

MACRO scs130lp_ebufn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ebufn_4 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.405 1.345 5.805 1.78 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.071 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.44 1.18 4.77 1.595 ;
        RECT 3.485 1.18 4.77 1.41 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.323 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.815 1.875 2.735 ;
        RECT 0.535 0.975 1.875 1.145 ;
        RECT 1.545 0.595 1.875 1.145 ;
        RECT 0.535 1.815 1.875 1.985 ;
        RECT 0.535 1.815 0.875 2.735 ;
        RECT 0.535 0.595 0.875 1.145 ;
        RECT 0.535 0.595 0.705 2.735 ;
        RECT 0.125 1.18 0.705 1.41 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.28 -0.085 5.61 1.135 ;
        RECT 3.265 -0.085 3.515 0.67 ;
        RECT 2.405 -0.085 2.735 0.965 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.21 2.525 5.54 3.415 ;
        RECT 3.545 2.865 3.875 3.415 ;
        RECT 2.545 2.695 2.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.71 1.95 6.145 3.075 ;
      RECT 5.975 0.255 6.145 3.075 ;
      RECT 4.325 2.185 6.145 2.355 ;
      RECT 2.045 2.015 4.495 2.185 ;
      RECT 2.045 1.475 2.215 2.185 ;
      RECT 0.875 1.475 2.215 1.645 ;
      RECT 0.875 1.315 1.885 1.645 ;
      RECT 5.78 0.255 6.145 1.135 ;
      RECT 4.665 1.765 5.11 2.015 ;
      RECT 4.94 0.255 5.11 2.015 ;
      RECT 4.195 0.34 5.11 1.01 ;
      RECT 4.78 0.255 5.11 1.01 ;
      RECT 4.085 2.525 4.415 3.075 ;
      RECT 3.045 2.355 3.375 3.075 ;
      RECT 0.115 2.905 2.375 3.075 ;
      RECT 2.045 2.355 2.375 3.075 ;
      RECT 1.045 2.155 1.375 3.075 ;
      RECT 0.115 1.815 0.365 3.075 ;
      RECT 3.045 2.525 4.415 2.695 ;
      RECT 2.045 2.355 3.375 2.525 ;
      RECT 2.055 1.135 3.085 1.305 ;
      RECT 2.915 0.255 3.085 1.305 ;
      RECT 2.055 0.255 2.225 1.305 ;
      RECT 2.915 0.84 4.025 1.01 ;
      RECT 3.695 0.255 4.025 1.01 ;
      RECT 0.115 0.255 0.365 1.01 ;
      RECT 1.045 0.255 1.375 0.805 ;
      RECT 0.115 0.255 2.225 0.425 ;
  END
END scs130lp_ebufn_4

MACRO scs130lp_ebufn_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ebufn_8 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.705 1.18 9.035 1.515 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.827 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.805 1.18 8.195 1.515 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.125 1.815 3.455 2.735 ;
        RECT 0.545 0.975 3.455 1.145 ;
        RECT 3.125 0.595 3.455 1.145 ;
        RECT 0.625 1.815 3.455 1.985 ;
        RECT 2.265 1.815 2.595 2.735 ;
        RECT 2.265 0.595 2.595 1.145 ;
        RECT 1.405 1.815 1.735 2.735 ;
        RECT 1.405 0.595 1.735 1.145 ;
        RECT 0.545 0.595 0.875 1.145 ;
        RECT 0.125 1.18 0.835 1.41 ;
        RECT 0.545 0.595 0.835 1.41 ;
        RECT 0.625 0.595 0.795 2.735 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 9.205 -0.085 9.455 1.095 ;
        RECT 8.345 -0.085 8.515 0.67 ;
        RECT 6.645 -0.085 6.815 0.965 ;
        RECT 5.785 -0.085 5.955 0.965 ;
        RECT 4.925 -0.085 5.095 0.965 ;
        RECT 3.985 -0.085 4.235 0.965 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 9.205 1.815 9.455 3.415 ;
        RECT 8.265 2.655 8.515 3.415 ;
        RECT 6.565 2.705 6.815 3.415 ;
        RECT 5.785 2.155 5.955 3.415 ;
        RECT 4.925 2.155 5.095 3.415 ;
        RECT 3.985 2.155 4.235 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.695 1.815 9.025 3.075 ;
      RECT 7.495 2.315 9.025 2.485 ;
      RECT 8.365 1.815 9.025 2.485 ;
      RECT 7.495 2.025 7.665 2.485 ;
      RECT 6.555 2.025 7.665 2.195 ;
      RECT 6.555 1.475 6.725 2.195 ;
      RECT 8.365 0.84 8.535 2.485 ;
      RECT 1.095 1.475 6.725 1.645 ;
      RECT 1.095 1.315 3.465 1.645 ;
      RECT 8.365 0.84 9.025 1.01 ;
      RECT 8.695 0.255 9.025 1.01 ;
      RECT 7.835 1.685 8.165 2.145 ;
      RECT 7.415 1.685 8.165 1.855 ;
      RECT 7.415 0.255 7.635 1.855 ;
      RECT 7.415 0.255 8.165 1.01 ;
      RECT 6.995 2.365 7.325 3.075 ;
      RECT 6.135 1.815 6.385 3.075 ;
      RECT 5.275 1.815 5.605 3.075 ;
      RECT 4.415 1.815 4.745 3.075 ;
      RECT 0.115 2.905 3.805 3.075 ;
      RECT 3.635 1.815 3.805 3.075 ;
      RECT 2.775 2.155 2.945 3.075 ;
      RECT 1.915 2.155 2.085 3.075 ;
      RECT 0.975 2.155 1.225 3.075 ;
      RECT 0.115 1.815 0.445 3.075 ;
      RECT 6.135 2.365 7.325 2.535 ;
      RECT 3.635 1.815 6.385 1.985 ;
      RECT 3.635 1.135 7.245 1.305 ;
      RECT 6.995 0.255 7.245 1.305 ;
      RECT 6.135 0.255 6.465 1.305 ;
      RECT 5.275 0.295 5.605 1.305 ;
      RECT 4.415 0.255 4.745 1.305 ;
      RECT 3.635 0.255 3.805 1.305 ;
      RECT 0.115 0.255 0.365 1.01 ;
      RECT 2.775 0.255 2.945 0.805 ;
      RECT 1.915 0.255 2.085 0.805 ;
      RECT 1.055 0.255 1.225 0.805 ;
      RECT 0.115 0.255 3.805 0.425 ;
  END
END scs130lp_ebufn_8

MACRO scs130lp_ebufn_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ebufn_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.49 1.245 0.835 2.15 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.507 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.44 1.175 3.77 1.78 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.405 1.175 2.755 2.89 ;
        RECT 1.905 1.005 2.575 1.175 ;
        RECT 2.12 2.025 2.45 3.075 ;
        RECT 1.905 0.595 2.405 1.175 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.085 -0.085 3.415 0.665 ;
        RECT 1.065 -0.085 1.395 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.94 1.815 3.27 3.415 ;
        RECT 1.345 2.395 1.675 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.875 1.985 4.205 2.665 ;
      RECT 4.035 0.255 4.205 2.665 ;
      RECT 1.21 1.185 1.735 1.515 ;
      RECT 1.565 0.255 1.735 1.515 ;
      RECT 2.745 0.835 4.205 1.005 ;
      RECT 3.875 0.255 4.205 1.005 ;
      RECT 2.745 0.255 2.915 1.005 ;
      RECT 1.565 0.255 2.915 0.425 ;
      RECT 0.125 2.395 0.455 3.075 ;
      RECT 0.125 2.395 1.175 2.565 ;
      RECT 1.005 1.685 1.175 2.565 ;
      RECT 0.125 0.635 0.295 3.075 ;
      RECT 1.005 1.685 2.235 1.855 ;
      RECT 1.905 1.345 2.235 1.855 ;
      RECT 0.125 0.635 0.485 1.075 ;
  END
END scs130lp_ebufn_lp

MACRO scs130lp_ebufn_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ebufn_lp2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 0.44 0.875 1.435 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.605 3.235 2.15 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.82 2.075 2.275 3.065 ;
        RECT 2.045 1.605 2.275 3.065 ;
        RECT 1.67 1.605 2.275 1.775 ;
        RECT 1.67 1.075 2 1.775 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.575 -0.085 2.905 1.075 ;
        RECT 1.055 -0.085 1.385 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.84 2.33 3.17 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.37 2.33 3.725 3.065 ;
      RECT 3.555 0.745 3.725 3.065 ;
      RECT 1.16 0.725 1.49 1.485 ;
      RECT 2.18 1.255 3.725 1.425 ;
      RECT 3.395 0.745 3.725 1.425 ;
      RECT 2.18 0.725 2.35 1.425 ;
      RECT 1.16 0.725 2.35 0.895 ;
      RECT 0.115 1.675 0.445 3.065 ;
      RECT 1.16 1.675 1.49 2.395 ;
      RECT 0.115 1.675 1.49 1.845 ;
      RECT 0.115 0.265 0.365 3.065 ;
  END
END scs130lp_ebufn_lp2

MACRO scs130lp_edfxbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_edfxbp_1 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.84 1.1 7.17 1.43 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.18 2.835 1.51 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 2.735 1.415 3.065 ;
        RECT 1.085 1.92 1.31 3.065 ;
    END
  END DE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5712 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.05 0.265 14.3 3.065 ;
        RECT 14.045 0.265 14.3 2.15 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5838 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.605 1.835 13.36 2.165 ;
        RECT 13.19 0.895 13.36 2.165 ;
        RECT 12.88 0.895 13.36 1.145 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 14.4 0.085 ;
        RECT 13.42 -0.085 13.75 0.365 ;
        RECT 12.37 -0.085 12.7 0.365 ;
        RECT 10.43 -0.085 10.76 0.365 ;
        RECT 7.7 -0.085 8.03 0.92 ;
        RECT 5.46 -0.085 5.79 0.895 ;
        RECT 1.565 -0.085 1.815 0.705 ;
        RECT 0.145 -0.085 0.395 1.335 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 14.4 3.415 ;
        RECT 13.54 2.695 13.87 3.415 ;
        RECT 12.56 2.695 12.89 3.415 ;
        RECT 10.87 2.785 11.04 3.415 ;
        RECT 7.72 2.31 7.89 3.415 ;
        RECT 5.98 2.065 6.23 3.415 ;
        RECT 1.92 2.095 2.09 3.415 ;
        RECT 0.145 2.385 0.395 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 12.095 1.92 12.385 2.15 ;
      RECT 3.455 1.92 3.745 2.15 ;
      RECT 3.455 1.965 12.385 2.105 ;
      RECT 8.255 1.55 8.545 1.78 ;
      RECT 4.895 1.55 5.185 1.78 ;
      RECT 4.895 1.595 8.545 1.735 ;
    LAYER li ;
      RECT 11.22 2.705 12.38 2.875 ;
      RECT 12.21 2.345 12.38 2.875 ;
      RECT 11.22 2.435 11.39 2.875 ;
      RECT 9.3 2.085 9.63 2.685 ;
      RECT 9.3 2.435 11.39 2.605 ;
      RECT 12.21 2.345 13.865 2.515 ;
      RECT 13.54 0.545 13.865 2.515 ;
      RECT 11.8 0.545 13.865 0.715 ;
      RECT 9.47 0.545 11.11 0.715 ;
      RECT 10.94 0.265 11.97 0.595 ;
      RECT 9.47 0.265 9.8 0.715 ;
      RECT 12.02 1.325 12.355 2.165 ;
      RECT 11.565 1.595 12.355 1.905 ;
      RECT 11.86 0.895 12.19 1.905 ;
      RECT 11.86 1.325 13.01 1.655 ;
      RECT 11.57 2.085 11.82 2.525 ;
      RECT 9.83 2.085 11.82 2.255 ;
      RECT 11.29 0.775 11.62 1.145 ;
      RECT 8.925 0.685 9.255 1.145 ;
      RECT 8.925 0.895 11.62 1.065 ;
      RECT 8.87 2.865 10.69 3.065 ;
      RECT 10.36 2.785 10.69 3.065 ;
      RECT 6.41 2.82 7.54 2.99 ;
      RECT 7.37 1.96 7.54 2.99 ;
      RECT 6.41 1.555 6.66 2.99 ;
      RECT 6.49 0.265 6.66 2.99 ;
      RECT 8.07 2.515 9.12 2.685 ;
      RECT 8.95 1.735 9.12 2.685 ;
      RECT 8.07 1.96 8.24 2.685 ;
      RECT 7.37 1.96 8.24 2.13 ;
      RECT 8.95 1.735 10.52 1.905 ;
      RECT 10.19 1.345 10.52 1.905 ;
      RECT 5.52 1.555 6.66 1.885 ;
      RECT 6.085 0.265 6.66 0.805 ;
      RECT 8.42 1.385 8.67 2.335 ;
      RECT 8.285 0.46 8.54 1.78 ;
      RECT 8.285 1.385 9.95 1.555 ;
      RECT 9.62 1.245 9.95 1.555 ;
      RECT 8.21 0.46 8.54 0.92 ;
      RECT 6.94 1.61 7.19 2.64 ;
      RECT 6.94 1.61 7.52 1.78 ;
      RECT 7.35 0.75 7.52 1.78 ;
      RECT 7.775 1.1 8.105 1.77 ;
      RECT 7.35 1.1 8.105 1.27 ;
      RECT 6.965 0.75 7.52 0.92 ;
      RECT 6.965 0.54 7.295 0.92 ;
      RECT 4.565 0.435 4.735 2.365 ;
      RECT 5.97 0.985 6.3 1.315 ;
      RECT 4.565 1.075 6.3 1.245 ;
      RECT 4.565 0.435 4.895 1.245 ;
      RECT 3.865 2.895 5.775 3.065 ;
      RECT 5.445 2.265 5.775 3.065 ;
      RECT 3.865 1.96 4.035 3.065 ;
      RECT 4.215 2.545 5.245 2.715 ;
      RECT 4.915 1.96 5.245 2.715 ;
      RECT 2.63 1.745 2.88 2.555 ;
      RECT 4.215 0.435 4.385 2.715 ;
      RECT 2.63 1.745 3.31 1.915 ;
      RECT 3.14 0.615 3.31 1.915 ;
      RECT 3.14 1.1 4.385 1.27 ;
      RECT 4.055 0.435 4.385 1.27 ;
      RECT 3.14 0.615 3.315 1.27 ;
      RECT 2.985 0.615 3.315 1 ;
      RECT 3.495 0.265 3.825 0.92 ;
      RECT 1.995 0.265 2.325 0.65 ;
      RECT 1.995 0.265 3.825 0.435 ;
      RECT 3.49 1.45 3.685 2.15 ;
      RECT 3.49 1.45 3.82 1.78 ;
      RECT 2.27 2.735 3.31 2.905 ;
      RECT 3.06 2.095 3.31 2.905 ;
      RECT 2.27 1.745 2.44 2.905 ;
      RECT 1.49 1.745 1.74 2.555 ;
      RECT 1.49 1.745 2.44 1.915 ;
      RECT 1.135 0.885 2.165 1.055 ;
      RECT 2.555 0.615 2.805 1 ;
      RECT 1.995 0.83 2.805 1 ;
      RECT 1.135 0.265 1.385 1.055 ;
      RECT 0.575 0.875 0.905 3.065 ;
      RECT 0.575 1.235 2.2 1.565 ;
      RECT 4.915 1.45 5.245 1.78 ;
  END
END scs130lp_edfxbp_1

MACRO scs130lp_einvn_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvn_0 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.21 1.375 2.975 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 1.21 0.875 2.215 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 0.685 1.835 3.055 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.6 0.775 1.365 1.04 ;
        RECT 1.195 -0.085 1.365 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.6 2.385 0.935 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.1 0.265 0.43 2.78 ;
      RECT 0.1 0.265 1.015 0.595 ;
  END
END scs130lp_einvn_0

MACRO scs130lp_einvn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvn_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.5 1.21 0.9 1.75 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.348 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.07 1.495 1.96 1.75 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.95 0.9 3.075 ;
        RECT 0.085 0.705 0.705 1.04 ;
        RECT 0.375 0.345 0.705 1.04 ;
        RECT 0.085 0.705 0.33 3.075 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.195 0.995 1.745 1.325 ;
        RECT 1.195 -0.085 1.61 1.325 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.195 1.92 1.63 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.8 1.92 2.315 2.565 ;
      RECT 2.13 0.265 2.315 2.565 ;
      RECT 1.915 0.265 2.315 1.27 ;
      RECT 1.78 0.265 2.315 0.63 ;
  END
END scs130lp_einvn_1

MACRO scs130lp_einvn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvn_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.195 3.275 1.525 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.537 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.55 0.84 0.945 1.51 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.903 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.975 1.705 3.265 3.075 ;
        RECT 2.11 1.705 3.265 1.875 ;
        RECT 2.495 0.595 2.835 0.885 ;
        RECT 2.495 0.595 2.735 1.875 ;
        RECT 2.11 1.705 2.37 2.155 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.645 -0.085 1.975 0.835 ;
        RECT 0.55 -0.085 0.88 0.56 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.505 2.665 1.835 3.415 ;
        RECT 0.6 2.02 0.93 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.215 1.005 2.325 1.175 ;
      RECT 2.145 0.255 2.325 1.175 ;
      RECT 3.005 0.255 3.265 1.025 ;
      RECT 1.215 0.255 1.475 1.175 ;
      RECT 2.145 0.255 3.265 0.425 ;
      RECT 2.505 2.325 2.805 3.075 ;
      RECT 2.54 2.045 2.805 3.075 ;
      RECT 1.1 2.02 1.335 3.075 ;
      RECT 1.1 2.325 2.805 2.495 ;
      RECT 1.1 2.02 1.405 2.495 ;
      RECT 0.1 1.68 0.43 2.485 ;
      RECT 0.1 1.68 1.94 1.85 ;
      RECT 1.77 1.345 1.94 1.85 ;
      RECT 0.1 0.355 0.37 2.485 ;
      RECT 1.77 1.345 2.1 1.535 ;
  END
END scs130lp_einvn_2

MACRO scs130lp_einvn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvn_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.425 1.765 1.75 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.071 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.47 1.745 4.725 2.86 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.512 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 0.595 2.245 1.5 ;
        RECT 1.845 1.92 2.175 2.735 ;
        RECT 1.945 0.595 2.175 2.735 ;
        RECT 0.825 1.075 2.245 1.245 ;
        RECT 1.845 0.595 2.245 1.245 ;
        RECT 0.905 1.92 2.175 2.09 ;
        RECT 0.905 1.92 1.235 2.735 ;
        RECT 0.825 0.595 1.155 1.245 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.895 -0.085 5.225 1.115 ;
        RECT 4.035 -0.085 4.365 0.885 ;
        RECT 3.175 -0.085 3.505 0.555 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.895 1.815 5.18 3.415 ;
        RECT 3.565 2.095 3.895 3.415 ;
        RECT 2.705 2.095 3.035 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.35 1.395 5.655 3.075 ;
      RECT 5.395 0.255 5.655 3.075 ;
      RECT 2.775 1.395 5.655 1.575 ;
      RECT 2.775 1.065 3.105 1.575 ;
      RECT 2.415 0.255 2.605 1.265 ;
      RECT 3.605 1.055 4.725 1.225 ;
      RECT 4.535 0.255 4.725 1.225 ;
      RECT 0.375 0.255 0.645 1.205 ;
      RECT 3.605 0.725 3.865 1.225 ;
      RECT 3.675 0.255 3.865 1.225 ;
      RECT 2.415 0.725 3.865 0.895 ;
      RECT 1.335 0.255 1.665 0.895 ;
      RECT 2.415 0.255 2.675 0.895 ;
      RECT 0.375 0.255 2.675 0.425 ;
      RECT 4.065 1.755 4.3 3.075 ;
      RECT 3.205 1.755 3.395 3.075 ;
      RECT 0.395 2.905 2.535 3.075 ;
      RECT 2.345 1.755 2.535 3.075 ;
      RECT 1.405 2.26 1.675 3.075 ;
      RECT 0.395 1.92 0.665 3.075 ;
      RECT 2.345 1.755 4.3 1.925 ;
  END
END scs130lp_einvn_4

MACRO scs130lp_einvn_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvn_8 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.355 1.185 6.135 1.515 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.827 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.21 0.775 1.645 ;
        RECT 0.105 1.21 0.415 2.96 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.935 1.665 8.265 2.735 ;
        RECT 6.305 1.14 8.225 1.875 ;
        RECT 8.005 0.595 8.225 2.735 ;
        RECT 7.075 1.14 7.405 2.735 ;
        RECT 7.145 0.595 7.335 2.735 ;
        RECT 6.215 1.685 6.545 2.735 ;
        RECT 6.305 0.69 6.475 2.735 ;
        RECT 5.355 0.69 6.475 1.015 ;
        RECT 5.355 1.685 8.265 1.875 ;
        RECT 5.355 1.685 5.685 2.735 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 4.53 -0.085 4.79 1.115 ;
        RECT 3.67 -0.085 3.93 1.115 ;
        RECT 2.81 -0.085 3.07 1.115 ;
        RECT 1.95 -0.085 2.21 1.115 ;
        RECT 0.095 -0.085 0.39 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 4.495 2.095 4.825 3.415 ;
        RECT 3.635 2.095 3.965 3.415 ;
        RECT 2.775 2.095 3.105 3.415 ;
        RECT 1.915 2.095 2.245 3.415 ;
        RECT 0.595 1.815 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.485 1.285 5.185 1.505 ;
      RECT 4.96 0.255 5.185 1.505 ;
      RECT 4.1 0.255 4.36 1.505 ;
      RECT 3.24 0.255 3.5 1.505 ;
      RECT 2.38 0.255 2.64 1.505 ;
      RECT 1.485 0.255 1.78 1.505 ;
      RECT 8.395 0.255 8.695 1.095 ;
      RECT 7.505 0.255 7.835 0.97 ;
      RECT 6.645 0.255 6.975 0.97 ;
      RECT 4.96 0.255 6.975 0.52 ;
      RECT 4.96 0.255 8.695 0.425 ;
      RECT 4.995 2.905 8.695 3.075 ;
      RECT 8.435 1.825 8.695 3.075 ;
      RECT 4.135 1.675 4.325 3.075 ;
      RECT 3.275 1.675 3.465 3.075 ;
      RECT 2.415 1.675 2.605 3.075 ;
      RECT 1.485 1.675 1.745 3.075 ;
      RECT 7.575 2.055 7.765 3.075 ;
      RECT 6.715 2.055 6.905 3.075 ;
      RECT 5.855 2.055 6.045 3.075 ;
      RECT 4.995 1.675 5.185 3.075 ;
      RECT 1.485 1.675 5.185 1.925 ;
      RECT 0.985 0.665 1.315 3.075 ;
      RECT 0.585 0.665 1.315 1.04 ;
      RECT 0.585 0.265 0.795 1.04 ;
  END
END scs130lp_einvn_8

MACRO scs130lp_einvn_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvn_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.44 2.275 0.67 ;
        RECT 1.78 0.3 2.11 0.67 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.58 0.935 2.15 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.725 1.18 2.275 3.065 ;
        RECT 1.725 0.85 2.2 3.065 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.91 -0.085 1.24 1.05 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.705 2.33 1.035 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.12 0.72 0.425 3.065 ;
      RECT 1.175 1.23 1.505 1.6 ;
      RECT 0.12 1.23 1.505 1.4 ;
      RECT 0.12 0.72 0.45 1.4 ;
  END
END scs130lp_einvn_lp

MACRO scs130lp_einvn_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvn_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.325 0.255 1.815 0.685 ;
    END
  END A
  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.33 0.805 0.685 ;
    END
  END TEB
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 0.855 1.825 2.925 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.695 0.855 1.155 1.185 ;
        RECT 0.985 -0.085 1.155 1.185 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.705 2.845 1.035 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.195 0.855 0.525 2.985 ;
      RECT 0.94 1.535 1.11 2.205 ;
      RECT 0.195 1.535 1.11 1.705 ;
  END
END scs130lp_einvn_m

MACRO scs130lp_einvp_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvp_0 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.84 1.835 2.12 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.56 0.84 0.925 1.75 ;
    END
  END TE
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2937 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 2.29 1.835 3.075 ;
        RECT 1.205 0.34 1.7 0.67 ;
        RECT 1.205 2.29 1.835 2.49 ;
        RECT 1.205 0.34 1.385 2.49 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.55 -0.085 0.88 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.62 2.43 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.12 1.93 0.45 3.015 ;
      RECT 0.12 1.93 1.035 2.26 ;
      RECT 0.12 0.395 0.38 3.015 ;
  END
END scs130lp_einvp_0

MACRO scs130lp_einvp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvp_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.455 1.79 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.18 1.825 1.515 ;
        RECT 1.045 1.18 1.825 1.39 ;
    END
  END TE
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5076 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.35 1.96 0.865 3.04 ;
        RECT 0.625 0.255 0.865 3.04 ;
        RECT 0.185 0.255 0.865 1.04 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.035 -0.085 1.825 1.01 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.16 2.035 1.53 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.7 1.685 2.03 2.425 ;
      RECT 1.035 1.685 2.275 1.865 ;
      RECT 1.995 0.7 2.275 1.865 ;
      RECT 1.035 1.56 1.415 1.865 ;
  END
END scs130lp_einvp_1

MACRO scs130lp_einvp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvp_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.995 1.21 3.255 1.75 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.411 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 2.665 0.74 3.065 ;
    END
  END TE
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.495 0.595 2.825 2.735 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.495 -0.085 1.825 0.895 ;
        RECT 0.54 -0.085 0.925 1.115 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.635 2.115 1.965 3.415 ;
        RECT 0.91 1.825 1.095 3.415 ;
        RECT 0.57 1.825 1.095 2.495 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.095 1.065 2.325 1.235 ;
      RECT 2.065 0.255 2.325 1.235 ;
      RECT 1.095 0.255 1.325 1.235 ;
      RECT 2.995 0.255 3.255 1.04 ;
      RECT 2.065 0.255 3.255 0.425 ;
      RECT 2.135 2.905 3.255 3.075 ;
      RECT 2.995 1.92 3.255 3.075 ;
      RECT 1.265 1.775 1.465 3.075 ;
      RECT 2.135 1.775 2.325 3.075 ;
      RECT 1.265 1.775 2.325 1.945 ;
      RECT 0.11 1.425 0.4 2.485 ;
      RECT 0.11 1.425 2.09 1.595 ;
      RECT 0.11 0.72 0.37 2.485 ;
  END
END scs130lp_einvp_2

MACRO scs130lp_einvp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvp_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.705 1.425 4.375 1.75 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.819 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.21 3.24 1.43 ;
        RECT 2.875 1.065 3.24 1.43 ;
    END
  END TE
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5204 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.545 1.385 5.665 1.555 ;
        RECT 5.365 0.325 5.665 1.555 ;
        RECT 4.935 1.385 5.225 2.735 ;
        RECT 3.965 1.92 5.225 2.09 ;
        RECT 4.545 1.385 5.225 2.09 ;
        RECT 4.545 0.615 4.795 2.09 ;
        RECT 3.455 1.085 4.795 1.255 ;
        RECT 4.465 0.615 4.795 1.255 ;
        RECT 3.965 1.92 4.265 2.735 ;
        RECT 3.455 0.605 3.785 1.255 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 2.285 -0.085 2.615 0.555 ;
        RECT 1.425 -0.085 1.755 0.7 ;
        RECT 0.6 -0.085 0.86 1.115 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 2.755 2.105 3.085 3.415 ;
        RECT 1.895 2.095 2.225 3.415 ;
        RECT 0.6 1.815 0.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.255 2.905 5.665 3.075 ;
      RECT 5.395 1.815 5.665 3.075 ;
      RECT 2.395 1.755 2.585 3.075 ;
      RECT 1.515 1.755 1.725 3.075 ;
      RECT 4.435 2.26 4.765 3.075 ;
      RECT 3.255 1.92 3.795 3.075 ;
      RECT 1.515 1.755 3.535 1.925 ;
      RECT 4.965 0.265 5.195 1.215 ;
      RECT 1.03 0.87 2.705 1.04 ;
      RECT 3.965 0.265 4.295 0.895 ;
      RECT 2.84 0.265 3.19 0.895 ;
      RECT 1.925 0.725 3.19 0.895 ;
      RECT 1.03 0.255 1.255 1.04 ;
      RECT 1.925 0.255 2.115 1.04 ;
      RECT 2.84 0.265 5.195 0.435 ;
      RECT 0.135 0.255 0.43 3.075 ;
      RECT 1.065 1.42 1.345 2.245 ;
      RECT 0.135 1.42 1.345 1.645 ;
  END
END scs130lp_einvp_4

MACRO scs130lp_einvp_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvp_8 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.295 1.345 7.985 1.595 ;
        RECT 6.295 1.21 7.245 1.595 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.323 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.805 1.75 ;
    END
  END TE
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.415 1.005 8.56 1.175 ;
        RECT 8.335 0.615 8.56 1.175 ;
        RECT 8.305 1.005 8.535 2.735 ;
        RECT 5.685 1.765 8.535 1.935 ;
        RECT 8.155 1.005 8.535 1.935 ;
        RECT 7.415 0.725 7.665 1.175 ;
        RECT 7.445 1.765 7.635 2.735 ;
        RECT 5.755 0.725 7.665 0.995 ;
        RECT 6.585 1.765 6.775 2.735 ;
        RECT 5.755 0.725 6.125 1.935 ;
        RECT 5.685 1.525 5.915 2.735 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 4.855 -0.085 5.085 1.04 ;
        RECT 3.965 -0.085 4.295 1.04 ;
        RECT 3.105 -0.085 3.435 1.04 ;
        RECT 2.245 -0.085 2.575 1.04 ;
        RECT 0.555 -0.085 0.855 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 4.83 1.89 5.09 3.415 ;
        RECT 3.97 1.89 4.225 3.415 ;
        RECT 3.105 1.89 3.37 3.415 ;
        RECT 2.245 1.89 2.505 3.415 ;
        RECT 0.455 1.92 0.725 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.815 1.21 5.585 1.38 ;
      RECT 5.255 0.275 5.585 1.38 ;
      RECT 4.465 0.255 4.685 1.38 ;
      RECT 3.605 0.255 3.795 1.38 ;
      RECT 2.745 0.255 2.935 1.38 ;
      RECT 1.815 0.255 2.075 1.38 ;
      RECT 8.73 0.275 9.025 1.095 ;
      RECT 7.835 0.275 8.165 0.825 ;
      RECT 5.255 0.275 8.165 0.555 ;
      RECT 5.255 0.275 9.025 0.445 ;
      RECT 5.26 2.905 8.995 3.075 ;
      RECT 8.705 1.815 8.995 3.075 ;
      RECT 4.395 1.55 4.66 3.075 ;
      RECT 3.54 1.55 3.8 3.075 ;
      RECT 2.675 1.55 2.935 3.075 ;
      RECT 1.785 1.55 2.075 3.075 ;
      RECT 7.805 2.105 8.135 3.075 ;
      RECT 6.945 2.105 7.275 3.075 ;
      RECT 6.085 2.105 6.415 3.075 ;
      RECT 5.26 1.55 5.515 3.075 ;
      RECT 1.785 1.55 5.515 1.72 ;
      RECT 0.945 1.93 1.615 3.075 ;
      RECT 0.945 1.855 1.315 3.075 ;
      RECT 1.025 0.255 1.315 3.075 ;
  END
END scs130lp_einvp_8

MACRO scs130lp_einvp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvp_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.44 0.835 0.67 ;
        RECT 0.34 0.265 0.67 0.67 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.439 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 0.44 1.795 1.41 ;
    END
  END TE
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.44845 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 0.85 0.465 3.065 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.035 -0.085 1.285 1.145 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.42 2.075 1.75 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.95 1.605 2.28 3.065 ;
      RECT 1.985 0.485 2.28 3.065 ;
      RECT 0.91 1.605 1.24 1.935 ;
      RECT 0.91 1.605 2.28 1.775 ;
  END
END scs130lp_einvp_lp

MACRO scs130lp_einvp_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_einvp_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.325 0.285 1.765 0.64 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.285 0.805 0.64 ;
    END
  END TE
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.47 0.82 1.8 2.925 ;
    END
  END Z
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.68 0.82 1.155 1.03 ;
        RECT 0.985 -0.085 1.155 1.03 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.74 2.785 0.95 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.17 1.535 0.52 2.985 ;
      RECT 0.855 1.535 1.025 2.205 ;
      RECT 0.17 1.535 1.025 1.705 ;
      RECT 0.17 0.835 0.5 2.985 ;
  END
END scs130lp_einvp_m

MACRO scs130lp_fa_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fa_0 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.87 1.57 2.95 1.82 ;
        RECT 0.87 1.57 1.12 2.025 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.01 1.755 6.575 2.125 ;
        RECT 6.125 1.19 6.575 2.125 ;
        RECT 3.13 1.755 6.575 1.925 ;
        RECT 1.4 1.99 3.3 2.32 ;
        RECT 3.13 1.755 3.3 2.32 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 1.365 5.835 1.585 ;
        RECT 5.505 1.295 5.835 1.585 ;
        RECT 1.69 1.23 3.79 1.4 ;
        RECT 3.45 1.13 3.79 1.585 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.625 0.495 0.955 ;
        RECT 0.085 2.5 0.425 3.075 ;
        RECT 0.085 0.625 0.325 3.075 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.305 1.405 7.595 2.945 ;
        RECT 7.345 0.35 7.595 2.945 ;
        RECT 7.155 0.35 7.595 0.68 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.69 -0.085 6.985 0.68 ;
        RECT 4.36 -0.085 4.69 0.855 ;
        RECT 3.45 -0.085 3.78 0.96 ;
        RECT 2.415 -0.085 2.745 0.72 ;
        RECT 0.665 -0.085 0.995 0.955 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.805 2.635 7.135 3.415 ;
        RECT 4.36 2.435 4.69 3.415 ;
        RECT 3.47 2.325 3.745 3.415 ;
        RECT 2.445 2.83 2.775 3.415 ;
        RECT 0.595 2.66 0.89 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.315 2.295 5.645 2.665 ;
      RECT 5.315 2.295 6.955 2.465 ;
      RECT 6.745 0.85 6.955 2.465 ;
      RECT 6.745 0.85 7.175 1.195 ;
      RECT 5.31 0.85 7.175 1.02 ;
      RECT 5.31 0.835 6.52 1.02 ;
      RECT 5.31 0.63 5.6 1.02 ;
      RECT 4.86 2.095 5.145 2.665 ;
      RECT 3.915 2.095 4.19 2.665 ;
      RECT 3.915 2.095 5.145 2.265 ;
      RECT 3.96 1.025 5.14 1.195 ;
      RECT 4.86 0.63 5.14 1.195 ;
      RECT 3.96 0.63 4.19 1.195 ;
      RECT 1.915 0.89 3.235 1.06 ;
      RECT 2.915 0.64 3.235 1.06 ;
      RECT 1.915 0.64 2.245 1.06 ;
      RECT 2.945 2.49 3.225 3.035 ;
      RECT 1.995 2.49 2.275 3.035 ;
      RECT 1.995 2.49 3.225 2.66 ;
      RECT 1.06 2.705 1.825 3.035 ;
      RECT 1.06 2.195 1.23 3.035 ;
      RECT 0.53 2.195 1.23 2.365 ;
      RECT 0.53 1.125 0.7 2.365 ;
      RECT 0.495 1.125 0.7 1.455 ;
      RECT 0.495 1.125 1.52 1.295 ;
      RECT 1.255 0.64 1.52 1.295 ;
      RECT 1.255 0.64 1.745 0.97 ;
  END
END scs130lp_fa_0

MACRO scs130lp_fa_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fa_1 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.915 1.185 6.63 1.825 ;
        RECT 3.45 1.185 6.63 1.355 ;
        RECT 3.45 1.165 5.495 1.355 ;
        RECT 3.45 1.095 3.935 1.355 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 1.865 3.715 2.94 ;
        RECT 3.365 1.865 3.715 2.12 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.815 0.375 3.075 ;
        RECT 0.085 0.255 0.365 3.075 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5733 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.795 1.815 8.075 3.075 ;
        RECT 7.84 0.255 8.075 3.075 ;
        RECT 7.64 0.255 8.075 1.02 ;
    END
  END SUM
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.504 LAYER met1 ;
      ANTENNAMAXAREACAR 2.253175 LAYER li ;
      ANTENNAMAXAREACAR 2.253175 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.865079 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.865079 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 6.815 1.92 7.105 2.15 ;
        RECT 1.055 1.965 7.105 2.105 ;
        RECT 2.495 1.92 2.785 2.15 ;
        RECT 1.055 1.92 1.345 2.15 ;
      LAYER li ;
        RECT 6.82 1.185 7.12 2.13 ;
        RECT 2.365 1.865 2.785 2.13 ;
        RECT 1.005 1.295 1.345 2.13 ;
    END
  END A
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.14 -0.085 7.47 0.675 ;
        RECT 4.515 -0.085 4.845 0.655 ;
        RECT 3.635 -0.085 3.935 0.795 ;
        RECT 2.56 -0.085 2.89 1.015 ;
        RECT 0.535 -0.085 1.2 1.045 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.285 2.64 7.615 3.415 ;
        RECT 4.845 2.205 5.035 3.415 ;
        RECT 4.705 2.205 5.035 2.47 ;
        RECT 3.885 2.1 4.12 3.415 ;
        RECT 2.57 2.64 2.9 3.415 ;
        RECT 0.555 2.64 0.885 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.605 2.3 7.625 2.47 ;
      RECT 7.29 1.19 7.625 2.47 ;
      RECT 5.605 2.1 5.875 2.47 ;
      RECT 7.29 1.19 7.66 1.52 ;
      RECT 7.29 0.845 7.47 2.47 ;
      RECT 5.665 0.845 7.47 1.015 ;
      RECT 5.665 0.665 6.97 1.015 ;
      RECT 1.63 2.3 1.92 2.655 ;
      RECT 1.7 0.73 1.92 2.655 ;
      RECT 0.555 2.3 1.92 2.47 ;
      RECT 0.555 1.215 0.795 2.47 ;
      RECT 1.7 1.525 5.7 1.695 ;
      RECT 0.535 1.215 0.795 1.545 ;
      RECT 1.7 0.73 1.985 1.695 ;
      RECT 4.105 0.825 5.495 0.995 ;
      RECT 5.015 0.385 5.495 0.995 ;
      RECT 4.105 0.465 4.345 0.995 ;
      RECT 5.205 1.865 5.435 2.43 ;
      RECT 4.29 1.865 4.535 2.43 ;
      RECT 4.29 1.865 5.435 2.035 ;
      RECT 3.08 2.3 3.335 2.66 ;
      RECT 2.09 2.3 2.39 2.66 ;
      RECT 2.09 2.3 3.335 2.47 ;
      RECT 2.155 1.185 3.28 1.355 ;
      RECT 3.06 0.73 3.28 1.355 ;
      RECT 2.155 0.73 2.39 1.355 ;
  END
END scs130lp_fa_1

MACRO scs130lp_fa_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fa_2 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.636 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.815 1.415 8.265 1.75 ;
        RECT 6.765 2.325 8.005 2.495 ;
        RECT 7.815 1.415 8.005 2.495 ;
        RECT 6.765 1.93 6.935 2.495 ;
        RECT 6.275 1.93 6.935 2.1 ;
        RECT 5.305 1.845 6.445 2.015 ;
        RECT 6.115 1.675 6.445 2.015 ;
        RECT 5.305 1.335 5.475 2.015 ;
        RECT 4.325 1.335 5.475 1.505 ;
        RECT 3.22 1.435 4.495 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.636 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.525 0.525 9.025 0.695 ;
        RECT 8.5 0.255 9.025 0.695 ;
        RECT 5.645 1.335 6.695 1.505 ;
        RECT 6.525 0.525 6.695 1.505 ;
        RECT 5.645 1.335 5.905 1.665 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.477 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.83 1.57 2.57 1.75 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.115 1.815 7.305 2.145 ;
        RECT 7.115 0.865 7.295 2.145 ;
        RECT 6.865 0.865 7.295 1.75 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.725 0.875 0.905 ;
        RECT 0.545 0.255 0.875 0.905 ;
        RECT 0.615 2.32 0.805 3.075 ;
        RECT 0.085 2.32 0.805 2.49 ;
        RECT 0.085 0.725 0.335 2.49 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 7.475 -0.085 7.805 0.355 ;
        RECT 6.455 -0.085 6.785 0.355 ;
        RECT 5.105 -0.085 5.81 0.825 ;
        RECT 3.165 -0.085 3.375 0.915 ;
        RECT 1.045 -0.085 1.325 0.71 ;
        RECT 0.115 -0.085 0.375 0.555 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 7.465 2.665 7.795 3.415 ;
        RECT 6.24 2.665 6.935 3.415 ;
        RECT 6.24 2.27 6.57 3.415 ;
        RECT 5.355 2.64 5.685 3.415 ;
        RECT 3.095 2.145 3.425 3.415 ;
        RECT 0.975 2.32 1.35 3.415 ;
        RECT 0.115 2.66 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 8.735 1.92 9.025 2.15 ;
      RECT 4.895 1.92 5.185 2.15 ;
      RECT 0.575 1.92 0.865 2.15 ;
      RECT 0.575 1.965 9.025 2.105 ;
    LAYER li ;
      RECT 8.68 0.865 9.025 2.495 ;
      RECT 7.465 1.075 7.645 1.545 ;
      RECT 7.465 1.075 9.025 1.245 ;
      RECT 4.705 0.995 6.18 1.165 ;
      RECT 5.98 0.705 6.18 1.165 ;
      RECT 4.705 0.64 4.935 1.165 ;
      RECT 4.795 2.29 5.125 2.89 ;
      RECT 5.855 2.2 6.07 2.87 ;
      RECT 4.795 2.29 6.07 2.47 ;
      RECT 5.81 2.2 6.07 2.47 ;
      RECT 4.245 2.075 4.505 2.745 ;
      RECT 3.605 2.075 4.505 2.245 ;
      RECT 3.605 1.785 3.775 2.245 ;
      RECT 2.87 1.785 3.775 1.955 ;
      RECT 2.87 1.085 3.04 1.955 ;
      RECT 0.855 1.425 1.66 1.595 ;
      RECT 1.49 1.23 1.66 1.595 ;
      RECT 1.49 1.23 3.04 1.4 ;
      RECT 3.545 0.64 3.715 1.255 ;
      RECT 2.87 1.085 3.715 1.255 ;
      RECT 3.545 0.64 4.535 0.97 ;
      RECT 2.665 0.37 2.995 0.915 ;
      RECT 1.635 0.37 1.965 0.71 ;
      RECT 1.635 0.37 2.995 0.54 ;
      RECT 1.52 2.82 2.915 2.99 ;
      RECT 2.585 2.145 2.915 2.99 ;
      RECT 1.52 2.32 1.85 2.99 ;
      RECT 2.02 1.92 2.28 2.64 ;
      RECT 0.505 1.92 2.28 2.15 ;
      RECT 0.505 1.075 0.685 2.15 ;
      RECT 0.505 1.075 1.225 1.245 ;
      RECT 1.055 0.88 1.225 1.245 ;
      RECT 1.055 0.88 2.475 1.05 ;
      RECT 2.145 0.71 2.475 1.05 ;
      RECT 4.675 1.675 5.125 2.12 ;
  END
END scs130lp_fa_2

MACRO scs130lp_fa_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fa_4 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.636 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.825 1.345 5.72 1.675 ;
        RECT 2.295 1.745 4.995 1.915 ;
        RECT 4.825 1.345 4.995 1.915 ;
        RECT 2.295 1.385 3.99 1.915 ;
        RECT 2.295 1.265 2.53 1.915 ;
        RECT 1.5 2.895 2.465 3.075 ;
        RECT 2.295 1.265 2.465 3.075 ;
        RECT 1.5 1.93 1.67 3.075 ;
        RECT 0.525 1.93 1.67 2.1 ;
        RECT 0.26 1.405 0.695 2.01 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.636 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.875 1.55 1.775 1.755 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.477 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.075 0.265 2.245 0.64 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.95 1.755 9.51 1.925 ;
        RECT 9.265 0.84 9.51 1.925 ;
        RECT 7.95 0.84 9.51 1.01 ;
        RECT 8.81 1.755 9 3.075 ;
        RECT 8.81 0.255 9 1.01 ;
        RECT 7.95 1.755 8.14 3.075 ;
        RECT 7.95 0.255 8.14 1.01 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.23 1.735 7.575 1.925 ;
        RECT 7.215 1.045 7.575 1.925 ;
        RECT 7.09 1.735 7.28 3.075 ;
        RECT 6.23 1.045 7.575 1.225 ;
        RECT 7.09 0.255 7.28 1.225 ;
        RECT 6.23 1.735 6.42 3.075 ;
        RECT 6.23 0.255 6.42 1.225 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 9.17 -0.085 9.5 0.67 ;
        RECT 8.31 -0.085 8.64 0.67 ;
        RECT 7.45 -0.085 7.78 0.875 ;
        RECT 6.59 -0.085 6.92 0.875 ;
        RECT 5.71 -0.085 6.04 0.53 ;
        RECT 3.445 -0.085 3.775 0.865 ;
        RECT 2.425 -0.085 2.755 1.04 ;
        RECT 0.575 -0.085 0.905 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 9.17 2.105 9.5 3.415 ;
        RECT 8.31 2.105 8.64 3.415 ;
        RECT 7.45 2.105 7.78 3.415 ;
        RECT 6.59 2.105 6.92 3.415 ;
        RECT 5.73 2.435 6.06 3.415 ;
        RECT 3.48 2.435 3.81 3.415 ;
        RECT 2.635 2.105 2.855 3.415 ;
        RECT 0.525 2.62 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 7.775 1.18 8.065 1.41 ;
      RECT 4.415 1.18 4.705 1.41 ;
      RECT 1.535 1.18 1.825 1.41 ;
      RECT 1.535 1.225 8.065 1.365 ;
    LAYER li ;
      RECT 4.43 2.095 4.745 2.765 ;
      RECT 4.43 2.095 6.06 2.265 ;
      RECT 5.89 0.7 6.06 2.265 ;
      RECT 5.89 1.395 7.045 1.565 ;
      RECT 4.495 0.7 6.06 1.03 ;
      RECT 4.2 1.385 4.655 1.575 ;
      RECT 4.475 1.2 4.655 1.575 ;
      RECT 3.98 2.095 4.26 2.765 ;
      RECT 3.025 2.095 3.275 2.765 ;
      RECT 3.025 2.095 4.26 2.265 ;
      RECT 3.055 1.045 4.235 1.215 ;
      RECT 4.025 0.765 4.235 1.215 ;
      RECT 3.055 0.765 3.265 1.215 ;
      RECT 1.84 2.055 2.115 2.725 ;
      RECT 1.945 1.21 2.115 2.725 ;
      RECT 1.595 0.81 1.945 1.38 ;
      RECT 0.205 1.065 1.415 1.235 ;
      RECT 1.085 0.81 1.415 1.235 ;
      RECT 0.205 0.705 0.405 1.235 ;
      RECT 0.095 2.18 0.345 2.85 ;
      RECT 1.11 2.28 1.32 2.61 ;
      RECT 0.095 2.28 1.32 2.45 ;
      RECT 0.095 2.18 0.355 2.45 ;
      RECT 7.745 1.18 9.095 1.515 ;
  END
END scs130lp_fa_4

MACRO scs130lp_fa_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fa_lp 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.365 0.44 7.235 0.67 ;
        RECT 6.905 0.265 7.235 0.67 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.04 2.165 9.135 2.335 ;
        RECT 8.82 1.605 9.135 2.335 ;
        RECT 4.435 1.18 4.71 1.565 ;
        RECT 3.125 1.235 4.71 1.405 ;
        RECT 3.605 2.1 4.21 2.27 ;
        RECT 3.605 1.235 3.775 2.27 ;
        RECT 3.125 1.235 3.775 1.565 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.939 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.39 1.815 8.61 1.985 ;
        RECT 8.28 1.605 8.61 1.985 ;
        RECT 6.8 1.55 7.08 1.985 ;
        RECT 3.955 1.75 4.56 1.92 ;
        RECT 3.955 1.59 4.225 1.92 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 0.405 0.545 0.865 ;
        RECT 0.115 0.405 0.445 2.935 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.115 2.075 10.47 3.065 ;
        RECT 10.3 0.31 10.47 3.065 ;
        RECT 10.115 0.31 10.47 1.04 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.27 -0.085 9.6 0.77 ;
        RECT 5.59 -0.085 5.92 0.935 ;
        RECT 4.49 -0.085 4.82 0.65 ;
        RECT 1.405 1.195 2.595 1.365 ;
        RECT 2.265 0.685 2.595 1.365 ;
        RECT 1.405 -0.085 1.575 1.365 ;
        RECT 1.005 -0.085 1.575 0.865 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.665 2.075 9.915 3.415 ;
        RECT 5.75 2.865 6.08 3.415 ;
        RECT 4.69 2.515 5.02 3.415 ;
        RECT 1.735 2.245 2.065 3.415 ;
        RECT 0.645 1.895 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.045 2.515 8.375 3.065 ;
      RECT 8.045 2.515 9.485 2.685 ;
      RECT 9.315 1.22 9.485 2.685 ;
      RECT 9.82 1.22 10.12 1.89 ;
      RECT 8.19 1.22 10.12 1.39 ;
      RECT 8.19 0.685 8.36 1.39 ;
      RECT 7.975 0.685 8.36 1.125 ;
      RECT 3.255 2.45 3.86 2.715 ;
      RECT 3.255 1.745 3.425 2.715 ;
      RECT 2.775 1.745 3.425 1.915 ;
      RECT 2.775 0.83 2.945 1.915 ;
      RECT 0.7 1.545 2.945 1.715 ;
      RECT 7.26 1.305 8.01 1.635 ;
      RECT 4.89 1.465 6.62 1.635 ;
      RECT 6.45 1.2 6.62 1.635 ;
      RECT 0.7 1.045 1.03 1.715 ;
      RECT 4.89 0.83 5.06 1.635 ;
      RECT 6.45 1.2 7.43 1.37 ;
      RECT 2.775 0.83 3.605 1.055 ;
      RECT 2.775 0.83 5.06 1 ;
      RECT 3.25 0.685 3.58 1.055 ;
      RECT 7.515 2.515 7.845 3.065 ;
      RECT 5.22 2.515 5.55 3.065 ;
      RECT 5.22 2.515 7.845 2.685 ;
      RECT 5.24 1.115 6.27 1.285 ;
      RECT 6.1 0.85 6.27 1.285 ;
      RECT 5.24 0.32 5.41 1.285 ;
      RECT 6.1 0.85 7.745 1.02 ;
      RECT 7.415 0.685 7.745 1.02 ;
      RECT 5.08 0.32 5.41 0.65 ;
      RECT 2.265 2.895 4.39 3.065 ;
      RECT 4.06 2.515 4.39 3.065 ;
      RECT 2.265 2.445 2.595 3.065 ;
      RECT 1.755 0.32 2.085 1.015 ;
      RECT 3.9 0.32 4.23 0.65 ;
      RECT 1.755 0.32 4.23 0.49 ;
      RECT 1.205 1.895 1.535 3.065 ;
      RECT 2.825 2.095 3.075 2.715 ;
      RECT 2.245 2.095 3.075 2.265 ;
      RECT 2.245 1.895 2.415 2.265 ;
      RECT 1.205 1.895 2.415 2.065 ;
  END
END scs130lp_fa_lp

MACRO scs130lp_fa_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fa_m 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.265 2.495 0.465 ;
        RECT 1.115 0.265 2.245 0.64 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.504 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.135 2.825 6.515 2.995 ;
        RECT 2.135 2.615 3.69 2.995 ;
        RECT 2.135 2.34 2.305 2.995 ;
        RECT 1.085 2.34 2.305 2.51 ;
        RECT 1.085 2.34 1.415 2.875 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 2.69 1.955 3.065 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.695 0.52 1.025 ;
        RECT 0.155 0.695 0.345 2.86 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.335 0.735 7.525 2.86 ;
        RECT 7.1 0.735 7.525 0.945 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.73 -0.085 6.92 0.905 ;
        RECT 4.62 -0.085 4.95 0.825 ;
        RECT 3.82 -0.085 4.03 0.905 ;
        RECT 2.515 0.645 2.845 0.835 ;
        RECT 2.675 -0.085 2.845 0.835 ;
        RECT 0.74 -0.085 0.93 0.935 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.83 2.125 7 3.415 ;
        RECT 3.87 2.425 7 2.595 ;
        RECT 6.67 2.125 7 2.595 ;
        RECT 4.68 2.065 4.89 2.595 ;
        RECT 2.485 2.265 4.04 2.435 ;
        RECT 3.82 2.065 4.04 2.435 ;
        RECT 2.485 2.065 2.815 2.435 ;
        RECT 0.525 2.005 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.58 1.915 5.965 2.245 ;
      RECT 5.795 0.705 5.965 2.245 ;
      RECT 6.985 1.125 7.155 1.795 ;
      RECT 5.795 1.125 7.155 1.295 ;
      RECT 5.58 0.705 5.965 1.035 ;
      RECT 1.53 0.835 1.74 2.145 ;
      RECT 0.525 1.365 5.615 1.535 ;
      RECT 1.47 0.835 1.8 1.535 ;
      RECT 0.525 1.205 0.695 1.535 ;
      RECT 4.25 1.005 5.32 1.175 ;
      RECT 5.13 0.705 5.32 1.175 ;
      RECT 4.25 0.705 4.44 1.175 ;
      RECT 5.11 1.715 5.32 2.245 ;
      RECT 4.25 1.715 4.46 2.245 ;
      RECT 4.25 1.715 5.32 1.885 ;
      RECT 1.98 1.015 3.265 1.185 ;
      RECT 3.055 0.735 3.265 1.185 ;
      RECT 1.98 0.835 2.31 1.185 ;
      RECT 1.96 1.715 2.17 2.145 ;
      RECT 3.055 1.715 3.265 2.085 ;
      RECT 1.96 1.715 3.265 1.885 ;
  END
END scs130lp_fa_m

MACRO scs130lp_fah_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fah_1 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.492 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.125 1.55 12.59 1.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.759 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.705 2.29 8.035 2.96 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.246 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.52 1.315 1.85 ;
    END
  END CI
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.975 2.895 2.585 3.065 ;
        RECT 2.335 2.68 2.585 3.065 ;
        RECT 1.515 0.44 2.09 0.67 ;
        RECT 1.76 0.28 2.09 0.67 ;
        RECT 0.635 0.74 1.685 0.91 ;
        RECT 1.515 0.44 1.685 0.91 ;
        RECT 0.975 2.03 1.145 3.065 ;
        RECT 0.635 2.03 1.145 2.2 ;
        RECT 0.635 0.74 0.805 2.2 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 0.44 0.445 3.065 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.44 0.085 ;
        RECT 12.645 -0.085 12.815 1.02 ;
        RECT 11.655 -0.085 11.905 0.67 ;
        RECT 7.615 -0.085 7.865 0.71 ;
        RECT 2.27 -0.085 2.44 0.67 ;
        RECT 0.66 -0.085 0.99 0.56 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.44 3.415 ;
        RECT 12.645 2.06 12.815 3.415 ;
        RECT 11.62 2.86 11.87 3.415 ;
        RECT 7.105 2.31 7.435 3.415 ;
        RECT 2.845 2.965 3.175 3.415 ;
        RECT 0.625 2.38 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 10.655 1.55 10.945 1.78 ;
      RECT 9.215 1.55 9.505 1.78 ;
      RECT 6.815 1.55 7.105 1.78 ;
      RECT 6.815 1.595 10.945 1.735 ;
      RECT 9.215 1.92 9.505 2.15 ;
      RECT 5.375 1.92 5.665 2.15 ;
      RECT 5.375 1.965 9.505 2.105 ;
      RECT 6.335 1.55 6.625 1.78 ;
      RECT 2.975 1.55 3.265 1.78 ;
      RECT 2.975 1.595 6.625 1.735 ;
    LAYER li ;
      RECT 12.995 0.34 13.325 3.065 ;
      RECT 11.445 1.2 11.775 1.675 ;
      RECT 11.445 1.2 13.325 1.37 ;
      RECT 12.135 2.06 12.465 3.065 ;
      RECT 8.335 2.875 10.07 3.045 ;
      RECT 9.74 2.68 10.07 3.045 ;
      RECT 8.335 1.24 8.505 3.045 ;
      RECT 9.74 2.68 11.44 2.85 ;
      RECT 11.27 2.51 12.465 2.68 ;
      RECT 8.335 1.24 8.71 1.41 ;
      RECT 8.54 0.265 8.71 1.41 ;
      RECT 9.785 0.265 10.115 1.08 ;
      RECT 11.305 0.85 12.465 1.02 ;
      RECT 12.135 0.34 12.465 1.02 ;
      RECT 11.305 0.265 11.475 1.02 ;
      RECT 8.54 0.265 11.475 0.435 ;
      RECT 8.685 1.59 9.015 2.695 ;
      RECT 8.685 2.33 11.09 2.5 ;
      RECT 10.76 1.96 11.09 2.5 ;
      RECT 10.76 1.96 11.265 2.13 ;
      RECT 11.095 1.2 11.265 2.13 ;
      RECT 8.89 0.615 9.06 1.76 ;
      RECT 10.875 0.615 11.125 1.37 ;
      RECT 10.25 1.61 10.58 2.15 ;
      RECT 10.25 1.61 10.915 1.78 ;
      RECT 10.685 1.55 10.915 1.78 ;
      RECT 9.195 1.94 9.92 2.15 ;
      RECT 9.75 1.26 9.92 2.15 ;
      RECT 9.75 1.26 10.5 1.43 ;
      RECT 10.33 0.615 10.5 1.43 ;
      RECT 10.33 0.615 10.66 1.255 ;
      RECT 6.755 1.96 6.925 3.065 ;
      RECT 6.755 1.96 7.435 2.13 ;
      RECT 7.265 0.265 7.435 2.13 ;
      RECT 7.265 0.89 8.36 1.06 ;
      RECT 8.045 0.39 8.36 1.06 ;
      RECT 4.37 0.265 7.435 0.435 ;
      RECT 3.355 2.895 6.575 3.065 ;
      RECT 6.405 1.96 6.575 3.065 ;
      RECT 4.705 2.68 5.68 3.065 ;
      RECT 3.355 2.615 3.525 3.065 ;
      RECT 2.765 2.615 3.525 2.785 ;
      RECT 1.325 2.075 1.665 2.715 ;
      RECT 1.495 1.09 1.665 2.715 ;
      RECT 4.705 1.81 4.875 3.065 ;
      RECT 2.765 2.33 2.935 2.785 ;
      RECT 1.325 2.33 2.935 2.5 ;
      RECT 6.045 1.96 6.575 2.13 ;
      RECT 4.16 1.81 4.875 1.98 ;
      RECT 6.045 1.055 6.215 2.13 ;
      RECT 4.16 1.35 4.33 1.98 ;
      RECT 3.815 1.35 4.33 1.68 ;
      RECT 1.17 1.09 1.665 1.34 ;
      RECT 5.34 1.055 6.215 1.225 ;
      RECT 5.34 0.965 5.67 1.225 ;
      RECT 5.895 2.33 6.225 2.715 ;
      RECT 5.055 2.33 6.225 2.5 ;
      RECT 5.055 1.405 5.225 2.5 ;
      RECT 2.375 1.2 2.705 1.58 ;
      RECT 4.99 0.965 5.16 1.575 ;
      RECT 2.375 1.2 3.14 1.37 ;
      RECT 2.97 0.615 3.14 1.37 ;
      RECT 4.91 0.965 5.16 1.295 ;
      RECT 3.67 0.965 5.16 1.135 ;
      RECT 3.67 0.615 3.84 1.135 ;
      RECT 2.97 0.615 3.84 0.785 ;
      RECT 4.195 2.16 4.525 2.715 ;
      RECT 3.115 2.265 4.525 2.435 ;
      RECT 3.115 1.98 3.285 2.435 ;
      RECT 1.865 1.98 3.285 2.15 ;
      RECT 1.865 0.85 2.195 2.15 ;
      RECT 1.865 0.85 2.79 1.02 ;
      RECT 2.62 0.265 2.79 1.02 ;
      RECT 5.885 0.615 6.215 0.875 ;
      RECT 4.02 0.615 6.215 0.785 ;
      RECT 4.02 0.265 4.19 0.785 ;
      RECT 2.62 0.265 4.19 0.435 ;
      RECT 3.465 1.915 3.98 2.085 ;
      RECT 3.465 1.61 3.635 2.085 ;
      RECT 3.32 0.965 3.49 1.78 ;
      RECT 3.005 1.55 3.49 1.78 ;
      RECT 9.24 0.615 9.57 1.76 ;
      RECT 6.755 0.665 7.085 1.78 ;
      RECT 6.395 0.615 6.575 1.78 ;
      RECT 5.405 1.405 5.865 2.15 ;
  END
END scs130lp_fah_1

MACRO scs130lp_fahcin_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fahcin_1 0 0 ;
  SIZE 12.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.46 1.345 0.805 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.759 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.66 1.18 5.155 1.67 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.561 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.245 1.08 8.575 1.41 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5644 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.365 0.44 7.555 0.885 ;
        RECT 6.525 1.96 6.855 2.715 ;
        RECT 6.525 0.295 6.695 2.715 ;
        RECT 6.365 0.295 6.695 0.885 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5922 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.12 0.375 12.37 3.065 ;
        RECT 11.825 0.375 12.37 1.075 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.48 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.48 0.085 ;
        RECT 11.315 -0.085 11.645 1.075 ;
        RECT 8.245 -0.085 8.575 0.9 ;
        RECT 5.225 -0.085 5.555 0.65 ;
        RECT 0.635 -0.085 0.805 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.48 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.48 3.415 ;
        RECT 11.69 1.855 11.94 3.415 ;
        RECT 8.495 1.94 8.665 3.415 ;
        RECT 5.145 2.785 5.475 3.415 ;
        RECT 0.555 2.055 0.885 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 10.175 1.55 10.465 1.78 ;
      RECT 6.815 1.55 7.105 1.78 ;
      RECT 3.935 1.55 4.225 1.78 ;
      RECT 1.535 1.55 1.825 1.78 ;
      RECT 1.535 1.595 10.465 1.735 ;
    LAYER li ;
      RECT 9.755 2.035 10.15 2.205 ;
      RECT 9.755 1.135 9.925 2.205 ;
      RECT 11.61 1.255 11.94 1.675 ;
      RECT 10.965 1.255 11.94 1.425 ;
      RECT 9.755 1.135 10.205 1.305 ;
      RECT 9.955 0.265 10.205 1.305 ;
      RECT 10.965 0.265 11.135 1.425 ;
      RECT 9.955 0.265 11.135 0.435 ;
      RECT 8.845 2.895 11.51 3.065 ;
      RECT 11.34 1.855 11.51 3.065 ;
      RECT 10.36 2.735 10.69 3.065 ;
      RECT 8.845 1.94 9.29 3.065 ;
      RECT 9.12 0.745 9.29 3.065 ;
      RECT 11.035 1.605 11.365 2.025 ;
      RECT 9.12 0.745 9.505 1.335 ;
      RECT 10.91 2.205 11.16 2.715 ;
      RECT 9.47 2.385 9.72 2.715 ;
      RECT 9.47 2.385 11.16 2.555 ;
      RECT 10.615 2.205 11.16 2.555 ;
      RECT 10.615 0.615 10.785 2.555 ;
      RECT 10.42 0.615 10.785 1.305 ;
      RECT 6.165 2.895 8.315 3.065 ;
      RECT 8.145 1.59 8.315 3.065 ;
      RECT 3.855 2.895 4.965 3.065 ;
      RECT 4.795 2.435 4.965 3.065 ;
      RECT 7.265 1.575 7.435 3.065 ;
      RECT 6.165 1.455 6.345 3.065 ;
      RECT 3.855 1.96 4.025 3.065 ;
      RECT 2.88 1.875 3.27 2.715 ;
      RECT 3.1 0.615 3.27 2.715 ;
      RECT 4.795 2.435 6.345 2.605 ;
      RECT 2.88 1.96 4.025 2.13 ;
      RECT 8.145 1.59 8.925 1.76 ;
      RECT 8.755 0.265 8.925 1.76 ;
      RECT 7.35 1.115 7.615 1.745 ;
      RECT 8.755 0.265 9.775 0.565 ;
      RECT 7.615 1.925 7.965 2.715 ;
      RECT 7.795 0.295 7.965 2.715 ;
      RECT 7.735 0.295 8.065 0.935 ;
      RECT 6.875 1.065 7.075 1.78 ;
      RECT 6.875 1.065 7.14 1.395 ;
      RECT 5.815 0.295 5.985 2.255 ;
      RECT 5.815 0.295 6.185 0.975 ;
      RECT 4.715 1.85 5.045 2.255 ;
      RECT 4.715 1.85 5.635 2.02 ;
      RECT 5.38 0.83 5.635 2.02 ;
      RECT 3.45 1.2 3.78 1.705 ;
      RECT 3.45 1.2 4.05 1.37 ;
      RECT 3.88 0.265 4.05 1.37 ;
      RECT 4.715 0.83 5.635 1 ;
      RECT 4.715 0.265 5.045 1 ;
      RECT 3.88 0.265 5.045 0.435 ;
      RECT 4.205 1.55 4.48 2.715 ;
      RECT 4.23 0.615 4.48 2.715 ;
      RECT 3.965 1.55 4.48 1.78 ;
      RECT 1.415 2.545 2.665 2.715 ;
      RECT 2.335 0.855 2.665 2.715 ;
      RECT 1.415 2.055 1.665 2.715 ;
      RECT 1.335 0.855 2.92 1.025 ;
      RECT 2.75 0.265 2.92 1.025 ;
      RECT 3.45 0.265 3.7 1.02 ;
      RECT 1.335 0.615 1.585 1.025 ;
      RECT 2.75 0.265 3.7 0.435 ;
      RECT 1.065 2.895 3.675 3.065 ;
      RECT 3.505 2.31 3.675 3.065 ;
      RECT 0.11 1.96 0.375 3.065 ;
      RECT 1.065 1.205 1.235 3.065 ;
      RECT 0.11 0.265 0.28 3.065 ;
      RECT 0.985 1.205 1.36 1.875 ;
      RECT 0.985 0.265 1.155 1.875 ;
      RECT 0.11 0.995 1.155 1.165 ;
      RECT 0.11 0.265 0.455 1.165 ;
      RECT 2.32 0.265 2.57 0.675 ;
      RECT 0.985 0.265 2.57 0.435 ;
      RECT 1.905 1.205 2.155 2.365 ;
      RECT 1.565 1.55 2.155 1.78 ;
      RECT 1.785 1.205 2.155 1.78 ;
      RECT 10.105 1.485 10.435 1.815 ;
  END
END scs130lp_fahcin_1

MACRO scs130lp_fahcon_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fahcon_1 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.345 0.805 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.005 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 1.18 5.05 1.53 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.561 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.705 1.18 8.035 1.515 ;
    END
  END CI
  PIN COUTN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0356 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.305 0.265 6.635 0.65 ;
        RECT 6.035 1.22 6.475 1.39 ;
        RECT 6.305 0.265 6.475 1.39 ;
        RECT 5.875 2.04 6.205 2.92 ;
        RECT 6.035 1.22 6.205 2.92 ;
    END
  END COUTN
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5796 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.155 0.265 11.42 3.065 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.52 0.085 ;
        RECT 10.61 -0.085 10.86 0.545 ;
        RECT 7.785 -0.085 8.035 1 ;
        RECT 4.845 -0.085 5.095 1 ;
        RECT 0.67 -0.085 0.84 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.52 3.415 ;
        RECT 10.66 2.285 10.91 3.415 ;
        RECT 7.32 1.86 7.65 3.415 ;
        RECT 4.565 1.775 4.895 3.415 ;
        RECT 0.655 1.96 0.985 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 9.215 0.81 9.505 1.04 ;
      RECT 6.815 0.81 7.105 1.04 ;
      RECT 5.855 0.81 6.145 1.04 ;
      RECT 2.015 0.81 2.305 1.04 ;
      RECT 2.015 0.855 9.505 0.995 ;
      RECT 8.735 1.92 9.025 2.15 ;
      RECT 6.335 1.92 6.625 2.15 ;
      RECT 2.975 1.92 3.265 2.15 ;
      RECT 2.975 1.965 9.025 2.105 ;
    LAYER li ;
      RECT 9.145 1.22 9.315 2.365 ;
      RECT 10.76 0.725 10.975 1.515 ;
      RECT 8.925 1.22 9.315 1.39 ;
      RECT 8.925 0.265 9.095 1.39 ;
      RECT 8.765 0.265 9.095 1.045 ;
      RECT 10.205 0.725 10.975 0.895 ;
      RECT 10.205 0.265 10.375 0.895 ;
      RECT 8.765 0.265 10.375 0.435 ;
      RECT 8.52 2.895 10.455 3.065 ;
      RECT 10.205 1.935 10.455 3.065 ;
      RECT 10.41 1.075 10.58 2.105 ;
      RECT 9.855 1.075 10.58 1.245 ;
      RECT 9.855 0.615 10.025 1.245 ;
      RECT 7.83 1.815 8.16 3.065 ;
      RECT 7.83 2.545 10.025 2.715 ;
      RECT 9.855 1.425 10.025 2.715 ;
      RECT 9.495 2.035 10.025 2.715 ;
      RECT 7.83 1.815 8.385 2.715 ;
      RECT 8.215 0.265 8.385 2.715 ;
      RECT 9.855 1.425 10.23 1.755 ;
      RECT 8.215 0.265 8.55 1.045 ;
      RECT 9.495 0.81 9.675 1.855 ;
      RECT 9.275 0.81 9.675 1.04 ;
      RECT 8.765 1.725 8.965 2.15 ;
      RECT 8.565 1.725 8.965 1.895 ;
      RECT 8.565 1.225 8.745 1.895 ;
      RECT 6.86 1.51 7.11 2.92 ;
      RECT 6.86 1.51 7.475 1.68 ;
      RECT 7.225 0.265 7.475 1.68 ;
      RECT 5.145 1.88 5.475 2.92 ;
      RECT 5.305 0.46 5.475 2.92 ;
      RECT 5.305 0.46 6.125 0.63 ;
      RECT 5.795 0.265 6.125 0.63 ;
      RECT 5.655 0.81 5.855 1.74 ;
      RECT 5.655 0.81 6.115 1.04 ;
      RECT 4.055 1.775 4.385 3.065 ;
      RECT 4.095 0.265 4.265 3.065 ;
      RECT 4.095 0.265 4.665 1 ;
      RECT 2.885 0.265 3.215 0.525 ;
      RECT 2.885 0.265 4.665 0.435 ;
      RECT 1.21 2.895 3.805 3.065 ;
      RECT 3.475 0.615 3.805 3.065 ;
      RECT 1.21 1.855 1.54 3.065 ;
      RECT 1.37 0.615 1.54 3.065 ;
      RECT 3.475 0.615 3.91 1.295 ;
      RECT 1.37 0.615 1.71 1.235 ;
      RECT 2.07 2.195 3.26 2.365 ;
      RECT 2.93 0.705 3.26 2.365 ;
      RECT 2.07 1.775 2.24 2.365 ;
      RECT 1.72 2.545 3.26 2.715 ;
      RECT 1.72 1.415 1.89 2.715 ;
      RECT 1.89 0.615 2.275 1.585 ;
      RECT 0.09 1.96 0.475 3.065 ;
      RECT 2.42 1.765 2.75 2.015 ;
      RECT 0.09 0.375 0.26 3.065 ;
      RECT 2.455 0.265 2.705 2.015 ;
      RECT 0.985 1.345 1.19 1.675 ;
      RECT 1.02 0.265 1.19 1.675 ;
      RECT 0.09 0.995 1.19 1.165 ;
      RECT 0.09 0.375 0.49 1.165 ;
      RECT 1.02 0.265 2.705 0.435 ;
      RECT 6.655 0.83 7.045 1.33 ;
      RECT 6.385 1.57 6.65 2.15 ;
  END
END scs130lp_fahcon_1

MACRO scs130lp_fill_1
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fill_1 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 0.48 0.085 ;
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 0.48 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_fill_1

MACRO scs130lp_fill_2
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fill_2 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_fill_2

MACRO scs130lp_fill_4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fill_4 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_fill_4

MACRO scs130lp_fill_8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_fill_8 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_fill_8

MACRO scs130lp_ha_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ha_0 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 1.055 2.8 1.385 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.915 3.27 2.295 ;
    END
  END B
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.255 2.435 4.715 3.075 ;
        RECT 4.435 0.375 4.715 3.075 ;
        RECT 4.355 0.375 4.715 1.425 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2937 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 2.495 0.5 3.075 ;
        RECT 0.095 0.385 0.425 1.425 ;
        RECT 0.095 0.385 0.325 3.075 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.855 -0.085 4.185 1.05 ;
        RECT 1.94 -0.085 2.27 0.545 ;
        RECT 0.595 -0.085 0.805 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.78 2.435 4.085 3.415 ;
        RECT 2.33 2.5 3.18 3.415 ;
        RECT 0.67 2.435 1 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.35 2.5 3.61 2.83 ;
      RECT 3.44 0.72 3.61 2.83 ;
      RECT 3.44 1.595 4.265 2.265 ;
      RECT 3.01 0.72 3.61 1.735 ;
      RECT 1.315 1.565 3.61 1.735 ;
      RECT 1.315 1.055 1.575 1.735 ;
      RECT 1.56 0.715 2.7 0.885 ;
      RECT 2.44 0.28 2.7 0.885 ;
      RECT 1.56 0.28 1.77 0.885 ;
      RECT 1.17 2.5 1.84 2.83 ;
      RECT 1.17 2.095 1.415 2.83 ;
      RECT 0.505 2.095 1.415 2.265 ;
      RECT 0.505 1.595 1.145 2.265 ;
      RECT 0.975 0.28 1.145 2.265 ;
      RECT 0.975 0.28 1.39 0.61 ;
  END
END scs130lp_ha_0

MACRO scs130lp_ha_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ha_1 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.315 1.57 2.79 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.96 1.23 3.27 1.76 ;
        RECT 1.885 1.23 3.27 1.4 ;
        RECT 1.885 1.18 2.145 1.85 ;
    END
  END B
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.395 0.29 4.715 3.075 ;
        RECT 4.325 0.29 4.715 1.09 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.74 0.505 3.075 ;
        RECT 0.095 0.26 0.365 3.075 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.79 -0.085 4.155 1.09 ;
        RECT 1.94 -0.085 2.27 0.67 ;
        RECT 0.535 -0.085 0.855 1.06 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.85 1.815 4.225 3.415 ;
        RECT 2.64 2.27 3.25 3.415 ;
        RECT 0.725 1.815 1.025 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.195 2.675 2.47 2.885 ;
      RECT 2.3 1.93 2.47 2.885 ;
      RECT 1.195 1.6 1.365 2.885 ;
      RECT 3.42 1.93 3.68 2.505 ;
      RECT 3.44 1.26 3.68 2.505 ;
      RECT 2.3 1.93 3.68 2.1 ;
      RECT 3.44 1.26 4.225 1.59 ;
      RECT 3.44 0.755 3.62 2.505 ;
      RECT 2.92 0.755 3.62 1.06 ;
      RECT 1.54 0.84 2.7 1.01 ;
      RECT 2.44 0.355 2.7 1.01 ;
      RECT 1.54 0.355 1.77 1.01 ;
      RECT 1.545 2.175 1.88 2.505 ;
      RECT 1.545 1.23 1.715 2.505 ;
      RECT 0.535 1.23 0.795 1.56 ;
      RECT 0.535 1.23 1.715 1.4 ;
      RECT 1.08 0.355 1.37 1.4 ;
  END
END scs130lp_ha_1

MACRO scs130lp_ha_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ha_2 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.495 0.815 1.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.495 1.315 1.795 ;
    END
  END B
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.45 0.255 3.725 2.305 ;
        RECT 3.39 0.255 3.725 1.015 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.31 1.695 4.645 3.075 ;
        RECT 4.465 0.255 4.645 3.075 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.825 -0.085 5.155 1.095 ;
        RECT 3.895 -0.085 4.225 1.015 ;
        RECT 2.795 -0.085 3.22 1.015 ;
        RECT 0.685 -0.085 0.935 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.815 1.815 5.015 3.415 ;
        RECT 3.81 2.815 4.14 3.415 ;
        RECT 2.95 2.815 3.28 3.415 ;
        RECT 1.78 2.255 1.995 3.415 ;
        RECT 0.32 1.975 0.65 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.165 2.475 4.14 2.645 ;
      RECT 3.97 1.185 4.14 2.645 ;
      RECT 1.11 1.965 1.39 2.635 ;
      RECT 2.165 1.685 2.335 2.645 ;
      RECT 1.11 1.965 1.655 2.135 ;
      RECT 1.485 0.65 1.655 2.135 ;
      RECT 1.485 1.685 2.335 1.855 ;
      RECT 1.485 0.65 1.66 1.855 ;
      RECT 3.97 1.185 4.295 1.515 ;
      RECT 1.485 0.65 1.805 0.98 ;
      RECT 2.505 1.185 2.695 2.305 ;
      RECT 1.84 1.185 3.28 1.515 ;
      RECT 1.84 1.15 2.335 1.515 ;
      RECT 1.975 0.7 2.335 1.515 ;
      RECT 0.185 1.075 1.315 1.245 ;
      RECT 1.105 0.65 1.315 1.245 ;
      RECT 0.185 0.65 0.515 1.245 ;
  END
END scs130lp_ha_2

MACRO scs130lp_ha_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ha_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.875 1.425 7.375 1.75 ;
        RECT 5.44 1.58 7.375 1.75 ;
        RECT 4.545 1.695 6.12 1.875 ;
        RECT 5.44 1.425 5.77 1.875 ;
        RECT 4.545 1.345 4.715 1.875 ;
        RECT 4.075 1.345 4.715 1.675 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.835 1.345 8.425 1.75 ;
        RECT 7.555 1.345 8.425 1.515 ;
        RECT 7.555 1.085 7.725 1.515 ;
        RECT 5.09 1.085 7.725 1.255 ;
        RECT 5.98 1.085 6.31 1.345 ;
        RECT 4.895 1.345 5.26 1.515 ;
        RECT 5.09 1.085 5.26 1.515 ;
    END
  END B
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.045 3.55 1.215 ;
        RECT 3.36 0.255 3.55 1.215 ;
        RECT 3.28 1.755 3.515 3.075 ;
        RECT 2.425 1.755 3.515 1.925 ;
        RECT 2.425 1.755 2.725 3.075 ;
        RECT 2.5 0.255 2.69 1.215 ;
        RECT 2.425 1.045 2.595 3.075 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.605 1.755 1.83 3.075 ;
        RECT 0.09 1.045 1.83 1.215 ;
        RECT 1.64 0.255 1.83 1.215 ;
        RECT 0.09 1.755 1.83 1.925 ;
        RECT 0.78 0.255 0.97 1.215 ;
        RECT 0.745 1.755 0.935 3.075 ;
        RECT 0.09 1.045 0.405 1.925 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.245 -0.085 8.445 0.755 ;
        RECT 7.83 -0.085 8.445 0.565 ;
        RECT 6.89 -0.085 7.22 0.535 ;
        RECT 5.605 -0.085 5.89 0.915 ;
        RECT 3.72 -0.085 4.06 0.805 ;
        RECT 2.86 -0.085 3.19 0.865 ;
        RECT 2 -0.085 2.33 0.67 ;
        RECT 1.14 -0.085 1.47 0.865 ;
        RECT 0.28 -0.085 0.61 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.95 2.63 9.52 3.415 ;
        RECT 9.295 2.105 9.52 3.415 ;
        RECT 7.34 2.95 7.685 3.415 ;
        RECT 5.56 2.385 5.89 3.415 ;
        RECT 4.68 2.385 5.01 3.415 ;
        RECT 3.685 2.195 4.015 3.415 ;
        RECT 2.895 2.095 3.11 3.415 ;
        RECT 2 1.81 2.255 3.415 ;
        RECT 1.105 2.095 1.435 3.415 ;
        RECT 0.245 2.095 0.575 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 9.215 0.81 9.505 1.04 ;
      RECT 2.015 0.81 2.305 1.04 ;
      RECT 2.015 0.855 9.505 0.995 ;
    LAYER li ;
      RECT 9.69 1.755 9.985 3.075 ;
      RECT 8.45 2.27 8.78 3.075 ;
      RECT 6.38 2.395 6.64 3.075 ;
      RECT 6.38 2.395 6.82 2.565 ;
      RECT 8.45 2.27 9.125 2.45 ;
      RECT 8.955 1.755 9.125 2.45 ;
      RECT 6.65 2.27 9.125 2.44 ;
      RECT 8.955 1.755 9.985 1.925 ;
      RECT 9.34 0.615 9.51 1.925 ;
      RECT 9.035 0.615 9.51 1.145 ;
      RECT 9.68 0.265 9.93 1.185 ;
      RECT 7.905 0.925 8.855 1.095 ;
      RECT 8.665 0.265 8.855 1.095 ;
      RECT 7.905 0.735 8.075 1.095 ;
      RECT 6.38 0.735 8.075 0.915 ;
      RECT 6.38 0.725 7.66 0.915 ;
      RECT 7.4 0.285 7.66 0.915 ;
      RECT 6.38 0.365 6.71 0.915 ;
      RECT 8.665 0.265 9.93 0.435 ;
      RECT 5.18 2.045 5.39 3.075 ;
      RECT 4.195 2.045 4.51 3.055 ;
      RECT 4.195 2.045 6.47 2.215 ;
      RECT 8.605 1.405 8.775 2.1 ;
      RECT 6.3 1.93 8.775 2.1 ;
      RECT 4.195 1.855 4.365 3.055 ;
      RECT 3.72 1.855 4.365 2.025 ;
      RECT 3.72 0.995 3.89 2.025 ;
      RECT 8.605 1.405 9.17 1.575 ;
      RECT 2.775 1.395 3.89 1.565 ;
      RECT 3.72 0.995 4.92 1.165 ;
      RECT 4.73 0.605 4.92 1.165 ;
      RECT 7.94 2.61 8.27 2.96 ;
      RECT 6.81 2.745 7.17 2.955 ;
      RECT 7 2.61 8.27 2.78 ;
      RECT 5.105 0.265 5.435 0.825 ;
      RECT 4.23 0.265 4.56 0.815 ;
      RECT 4.23 0.265 5.435 0.435 ;
      RECT 0.675 1.395 2.245 1.565 ;
      RECT 2.075 0.84 2.245 1.565 ;
  END
END scs130lp_ha_4

MACRO scs130lp_ha_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ha_lp 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.785 1.45 3.205 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.215 1.96 3.685 2.13 ;
        RECT 3.385 1.605 3.685 2.13 ;
        RECT 2.215 1.96 2.755 2.89 ;
        RECT 2.215 1.605 2.545 2.89 ;
    END
  END B
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.745 2.075 5.17 3.065 ;
        RECT 4.925 0.44 5.17 3.065 ;
        RECT 4.84 0.44 5.17 1.045 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.11 2.865 0.975 3.035 ;
        RECT 0.645 2.155 0.975 3.035 ;
        RECT 0.11 0.44 0.44 3.035 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.05 -0.085 4.38 1.045 ;
        RECT 2.25 -0.085 2.58 0.57 ;
        RECT 0.9 -0.085 1.15 1.335 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.215 2.075 4.545 3.415 ;
        RECT 3.01 2.31 3.34 3.415 ;
        RECT 1.175 2.075 1.505 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.59 2.31 4.035 3.065 ;
      RECT 3.865 1.225 4.035 3.065 ;
      RECT 4.355 1.225 4.685 1.895 ;
      RECT 1.68 1.1 1.985 1.43 ;
      RECT 3.42 1.225 4.685 1.395 ;
      RECT 3.26 0.605 3.59 1.27 ;
      RECT 1.68 1.1 3.59 1.27 ;
      RECT 1.82 0.75 3.01 0.92 ;
      RECT 2.76 0.265 3.01 0.92 ;
      RECT 1.82 0.265 2.07 0.92 ;
      RECT 1.705 1.725 2.035 3.065 ;
      RECT 0.87 1.725 2.035 1.895 ;
      RECT 0.87 1.565 1.5 1.895 ;
      RECT 1.33 0.265 1.5 1.895 ;
      RECT 1.33 0.265 1.64 0.645 ;
  END
END scs130lp_ha_lp

MACRO scs130lp_ha_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_ha_m 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.05 2.43 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 1.91 3.29 2.12 ;
        RECT 2.96 1.295 3.29 2.12 ;
    END
  END B
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.425 0.47 4.645 2.86 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 2.49 1.09 2.86 ;
        RECT 0.095 0.47 0.425 2.86 ;
    END
  END SUM
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.995 -0.085 4.185 0.935 ;
        RECT 1.99 -0.085 2.32 0.415 ;
        RECT 0.605 -0.085 0.795 0.74 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.995 2.125 4.185 3.415 ;
        RECT 2.79 2.49 3.12 3.415 ;
        RECT 1.27 2.43 1.48 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.47 0.795 3.8 3.025 ;
      RECT 1.325 1.56 2.78 1.73 ;
      RECT 2.61 0.945 2.78 1.73 ;
      RECT 1.325 1.06 1.495 1.73 ;
      RECT 2.61 0.945 3.8 1.115 ;
      RECT 3.05 0.795 3.8 1.115 ;
      RECT 1.54 0.595 2.77 0.765 ;
      RECT 2.56 0.345 2.77 0.765 ;
      RECT 1.54 0.345 1.75 0.765 ;
      RECT 1.68 2.36 2.125 2.57 ;
      RECT 1.68 1.95 1.85 2.57 ;
      RECT 0.605 1.95 1.85 2.12 ;
      RECT 0.975 0.345 1.145 2.12 ;
      RECT 0.605 1.45 0.775 2.12 ;
      RECT 0.975 0.345 1.3 0.675 ;
  END
END scs130lp_ha_m

MACRO scs130lp_inputiso0n_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inputiso0n_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.345 1.395 1.09 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.855 0.465 3.275 3.075 ;
    END
  END X
  PIN sleepb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.315 1.395 1.985 1.75 ;
    END
  END sleepb
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.44 -0.085 2.335 0.84 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.99 2.295 2.675 3.415 ;
        RECT 0.29 2.49 0.62 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.08 1.955 1.41 2.82 ;
      RECT 1.08 1.955 2.685 2.125 ;
      RECT 2.275 1.055 2.685 2.125 ;
      RECT 0.65 1.055 2.685 1.225 ;
      RECT 0.65 0.51 0.98 1.225 ;
  END
END scs130lp_inputiso0n_lp

MACRO scs130lp_inputiso0p_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inputiso0p_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 1.395 2.65 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.4 0.465 3.755 3.075 ;
    END
  END X
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 1.16 0.92 1.895 ;
    END
  END sleep
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.55 -0.085 2.885 0.835 ;
        RECT 0.895 -0.085 1.575 0.84 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.525 2.295 2.91 3.415 ;
        RECT 0.895 2.445 1.225 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.765 1.955 1.975 2.855 ;
      RECT 1.765 1.955 3.23 2.125 ;
      RECT 2.82 1.005 3.23 2.125 ;
      RECT 2.095 1.005 3.23 1.225 ;
      RECT 2.095 0.43 2.305 1.225 ;
      RECT 0.155 0.43 0.375 2.855 ;
      RECT 0.155 2.065 1.595 2.235 ;
      RECT 1.2 1.39 1.595 2.235 ;
  END
END scs130lp_inputiso0p_lp

MACRO scs130lp_inputiso1n_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inputiso1n_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.91 1.395 2.58 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.395 0.465 3.755 3.075 ;
    END
  END X
  PIN sleepb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.54 1.16 1.16 1.99 ;
    END
  END sleepb
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.525 -0.085 2.855 0.885 ;
        RECT 0.885 -0.085 1.215 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.525 2.295 2.91 3.415 ;
        RECT 1.19 2.5 1.52 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.095 1.955 2.305 2.88 ;
      RECT 2.095 1.955 3.225 2.125 ;
      RECT 2.895 1.055 3.225 2.125 ;
      RECT 1.87 1.055 3.225 1.225 ;
      RECT 1.87 0.43 2.065 1.225 ;
      RECT 1.735 0.43 2.065 0.885 ;
      RECT 0.345 2.16 0.59 2.82 ;
      RECT 0.125 2.16 1.7 2.33 ;
      RECT 1.37 1.315 1.7 2.33 ;
      RECT 0.125 0.885 0.37 2.33 ;
      RECT 0.12 0.43 0.365 0.885 ;
  END
END scs130lp_inputiso1n_lp

MACRO scs130lp_inputiso1p_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inputiso1p_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 1.35 1.225 1.75 ;
        RECT 0.555 1.16 0.855 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.855 0.465 3.275 3.075 ;
    END
  END X
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.435 1.35 2.105 1.75 ;
    END
  END sleep
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.01 -0.085 2.34 0.84 ;
        RECT 0.46 -0.085 0.76 0.84 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.56 2.295 2.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.77 1.955 1.1 2.82 ;
      RECT 0.77 1.955 2.685 2.125 ;
      RECT 2.35 1.01 2.685 2.125 ;
      RECT 1.28 1.01 2.685 1.18 ;
      RECT 1.28 0.44 1.49 1.18 ;
  END
END scs130lp_inputiso1p_lp

MACRO scs130lp_inputisolatch_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inputisolatch_lp 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.255 0.835 1.78 ;
        RECT 0.125 2.185 0.585 2.515 ;
        RECT 0.125 1.255 0.295 2.515 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4597 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.45 0.44 7.085 2.955 ;
    END
  END Q
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.355 1.45 4.685 1.78 ;
    END
  END SLEEPB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 5.95 -0.085 6.28 1.325 ;
        RECT 4.6 -0.085 4.85 0.905 ;
        RECT 2.97 -0.085 3.22 0.775 ;
        RECT 0.59 -0.085 0.92 0.745 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 5.865 1.915 6.195 3.415 ;
        RECT 4.775 2.29 5.155 3.415 ;
        RECT 2.515 2.125 2.845 3.415 ;
        RECT 0.13 2.685 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.515 2.905 4.605 3.075 ;
      RECT 4.435 1.95 4.605 3.075 ;
      RECT 5.335 1.915 5.665 2.955 ;
      RECT 5.495 0.445 5.665 2.955 ;
      RECT 3.515 1.785 3.845 3.075 ;
      RECT 4.435 1.95 5.665 2.12 ;
      RECT 5.46 0.445 5.665 0.775 ;
      RECT 1.495 2.29 1.855 2.735 ;
      RECT 1.685 1.33 1.855 2.735 ;
      RECT 4.895 1.075 5.225 1.745 ;
      RECT 1.575 0.345 1.745 1.5 ;
      RECT 4.15 1.075 5.225 1.245 ;
      RECT 2.415 0.945 3.56 1.115 ;
      RECT 3.39 0.255 3.56 1.115 ;
      RECT 4.15 0.255 4.32 1.245 ;
      RECT 2.415 0.555 2.585 1.115 ;
      RECT 1.575 0.555 2.585 0.725 ;
      RECT 1.575 0.345 1.97 0.725 ;
      RECT 3.39 0.255 4.32 0.425 ;
      RECT 4.015 2.055 4.265 2.735 ;
      RECT 4.015 1.445 4.185 2.735 ;
      RECT 2.075 1.445 4.185 1.615 ;
      RECT 2.075 1.285 3.98 1.615 ;
      RECT 3.73 0.595 3.98 1.615 ;
      RECT 2.075 0.895 2.245 1.615 ;
      RECT 1.915 0.895 2.245 1.16 ;
      RECT 3.045 1.785 3.295 3.075 ;
      RECT 1.155 2.905 2.345 3.075 ;
      RECT 2.175 1.785 2.345 3.075 ;
      RECT 1.155 1.95 1.325 3.075 ;
      RECT 1.185 1.67 1.515 2.12 ;
      RECT 2.175 1.785 3.295 1.955 ;
      RECT 1.185 0.915 1.355 2.12 ;
      RECT 0.16 0.915 1.355 1.085 ;
      RECT 0.16 0.345 0.41 1.085 ;
  END
END scs130lp_inputisolatch_lp

MACRO scs130lp_inv_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_0 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.955 0.4 2.12 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 0.395 0.875 2.97 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
        RECT 0.105 -0.085 0.4 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
        RECT 0.105 2.29 0.4 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_0

MACRO scs130lp_inv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_1 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.435 1.75 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 0.255 0.875 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
        RECT 0.105 -0.085 0.435 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
        RECT 0.105 1.92 0.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_1

MACRO scs130lp_inv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_16 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 5.04 LAYER li ;
      ANTENNAGATEAREA 5.04 LAYER met1 ;
      ANTENNAMAXAREACAR 0.021409 LAYER li ;
      ANTENNAMAXAREACAR 0.021409 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.026786 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.026786 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.005734 LAYER mcon ;
    PORT
      LAYER li ;
        RECT 6.225 1.335 6.485 1.75 ;
        RECT 5.365 1.335 5.625 1.75 ;
        RECT 4.505 1.335 4.765 1.75 ;
        RECT 3.645 1.335 3.905 1.75 ;
        RECT 2.785 1.335 3.045 1.75 ;
        RECT 1.925 1.335 2.185 1.75 ;
        RECT 1.065 1.335 1.325 1.75 ;
      LAYER met1 ;
        RECT 1.05 1.55 6.5 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    ANTENNADIFFAREA 4.704 LAYER met1 ;
    PORT
      LAYER li ;
        RECT 6.655 0.305 6.915 3.05 ;
        RECT 5.795 0.305 6.055 3.05 ;
        RECT 4.935 0.305 5.195 3.05 ;
        RECT 4.075 0.305 4.335 3.05 ;
        RECT 3.215 0.305 3.475 3.05 ;
        RECT 2.355 0.305 2.615 3.05 ;
        RECT 1.495 0.305 1.755 3.05 ;
        RECT 0.635 0.305 0.895 3.05 ;
      LAYER met1 ;
        RECT 0.62 1.92 6.93 2.15 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.085 -0.085 7.38 1.005 ;
        RECT 6.225 -0.085 6.485 1.005 ;
        RECT 5.365 -0.085 5.625 1.005 ;
        RECT 4.505 -0.085 4.765 1.005 ;
        RECT 3.645 -0.085 3.905 1.005 ;
        RECT 2.785 -0.085 3.045 1.005 ;
        RECT 1.925 -0.085 2.185 1.005 ;
        RECT 1.065 -0.085 1.325 1.005 ;
        RECT 0.17 -0.085 0.465 1.005 ;
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.085 1.92 7.38 3.415 ;
        RECT 6.225 1.92 6.485 3.415 ;
        RECT 5.365 1.92 5.625 3.415 ;
        RECT 4.505 1.92 4.765 3.415 ;
        RECT 3.645 1.92 3.905 3.415 ;
        RECT 2.785 1.92 3.045 3.415 ;
        RECT 1.925 1.92 2.185 3.415 ;
        RECT 1.065 1.92 1.325 3.415 ;
        RECT 0.17 1.92 0.465 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_16

MACRO scs130lp_inv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_2 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.435 1.75 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 0.305 0.835 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 1.005 -0.085 1.295 1.205 ;
        RECT 0.105 -0.085 0.435 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 1.005 1.815 1.295 3.415 ;
        RECT 0.105 1.92 0.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_2

MACRO scs130lp_inv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_4 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.21 1.845 1.515 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.56 1.755 2.3 1.925 ;
        RECT 2.025 0.84 2.3 1.925 ;
        RECT 0.565 0.87 2.3 1.04 ;
        RECT 1.425 0.84 2.3 1.04 ;
        RECT 1.42 1.755 1.685 3.075 ;
        RECT 1.425 0.255 1.685 1.04 ;
        RECT 0.56 1.755 0.825 3.075 ;
        RECT 0.565 0.255 0.825 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.855 -0.085 2.15 0.67 ;
        RECT 0.995 -0.085 1.255 0.7 ;
        RECT 0.1 -0.085 0.395 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.855 2.095 2.15 3.415 ;
        RECT 0.995 2.095 1.25 3.415 ;
        RECT 0.1 1.815 0.39 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_4

MACRO scs130lp_inv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_8 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.425 1.395 3.815 1.585 ;
        RECT 2.06 1.385 3.815 1.585 ;
        RECT 2.06 1.16 2.365 1.585 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.755 4.225 1.925 ;
        RECT 3.985 1.045 4.225 1.925 ;
        RECT 2.535 1.045 4.225 1.215 ;
        RECT 3.395 1.755 3.655 3.075 ;
        RECT 3.395 0.255 3.655 1.215 ;
        RECT 2.535 1.755 2.795 3.075 ;
        RECT 2.535 0.255 2.795 1.215 ;
        RECT 1.675 0.82 2.795 0.99 ;
        RECT 1.675 1.755 1.935 3.075 ;
        RECT 1.675 0.255 1.935 0.99 ;
        RECT 0.085 1.045 1.89 1.215 ;
        RECT 1.675 0.255 1.89 1.215 ;
        RECT 0.815 1.755 1.075 3.075 ;
        RECT 0.815 0.255 1.075 1.215 ;
        RECT 0.085 1.045 0.255 1.925 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.825 -0.085 4.12 0.875 ;
        RECT 2.965 -0.085 3.225 0.875 ;
        RECT 2.105 -0.085 2.365 0.65 ;
        RECT 1.245 -0.085 1.505 0.875 ;
        RECT 0.35 -0.085 0.645 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.825 2.095 4.12 3.415 ;
        RECT 2.965 2.095 3.225 3.415 ;
        RECT 2.105 2.095 2.365 3.415 ;
        RECT 1.245 2.095 1.505 3.415 ;
        RECT 0.35 2.105 0.645 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_8

MACRO scs130lp_inv_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_lp 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.955 0.835 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.96 1.315 3 ;
        RECT 1.085 0.315 1.315 3 ;
        RECT 0.985 0.315 1.315 0.775 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.165 -0.085 0.495 0.775 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.455 1.96 0.785 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_lp

MACRO scs130lp_inv_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_inv_m 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.955 0.355 2.12 ;
        RECT 0.155 0.84 0.325 2.12 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 0.445 0.805 2.96 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
        RECT 0.165 -0.085 0.355 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
        RECT 0.165 2.3 0.375 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_inv_m

MACRO scs130lp_invkapwr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invkapwr_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.79 0.475 1.8 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.645 0.84 1.285 1.9 ;
        RECT 0.645 0.84 0.875 2.88 ;
        RECT 0.645 0.395 0.845 2.88 ;
    END
  END Y
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 1.37 2.945 ;
      LAYER li ;
        RECT 1.045 2.18 1.345 2.945 ;
        RECT 0.155 2.18 0.475 2.945 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 1.015 -0.085 1.345 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_invkapwr_1

MACRO scs130lp_invkapwr_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invkapwr_2 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.693 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.415 1.21 1.425 1.545 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8043 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.715 1.78 1.885 ;
        RECT 1.595 0.84 1.78 1.885 ;
        RECT 1.1 0.84 1.78 1.04 ;
        RECT 1.1 0.395 1.325 1.04 ;
        RECT 1.01 1.715 1.27 3.045 ;
        RECT 0.155 1.715 0.41 3.045 ;
    END
  END Y
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 1.85 2.945 ;
      LAYER li ;
        RECT 1.44 2.055 1.695 3.075 ;
        RECT 0.58 2.055 0.84 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.495 -0.085 1.825 0.67 ;
        RECT 0.635 -0.085 0.93 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_invkapwr_2

MACRO scs130lp_invkapwr_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invkapwr_4 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.386 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 1.21 2.865 1.545 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.23 1.715 3.22 1.885 ;
        RECT 3.035 0.84 3.22 1.885 ;
        RECT 0.23 0.84 3.22 1.04 ;
        RECT 2.45 1.715 2.71 3.045 ;
        RECT 2.02 0.395 2.275 1.04 ;
        RECT 1.595 1.715 1.85 3.045 ;
        RECT 1.16 0.395 1.42 1.04 ;
        RECT 0.735 1.715 0.99 3.045 ;
        RECT 0.23 0.84 0.4 1.885 ;
    END
  END Y
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 3.29 2.945 ;
      LAYER li ;
        RECT 2.88 2.055 3.135 3.075 ;
        RECT 2.02 2.055 2.28 3.075 ;
        RECT 1.16 2.055 1.42 3.075 ;
        RECT 0.3 2.055 0.56 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.445 -0.085 2.745 0.67 ;
        RECT 1.59 -0.085 1.85 0.67 ;
        RECT 0.695 -0.085 0.99 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_invkapwr_4

MACRO scs130lp_invkapwr_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invkapwr_8 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.772 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.515 1.21 5.265 1.54 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.175 1.71 5.62 1.885 ;
        RECT 5.435 0.84 5.62 1.885 ;
        RECT 0.175 0.84 5.62 1.04 ;
        RECT 4.93 1.71 5.19 3.045 ;
        RECT 4.075 1.71 4.33 3.045 ;
        RECT 4.07 0.395 4.33 1.04 ;
        RECT 3.215 1.71 3.47 3.045 ;
        RECT 3.21 0.395 3.47 1.04 ;
        RECT 2.355 1.71 2.61 3.045 ;
        RECT 2.35 0.395 2.61 1.04 ;
        RECT 1.495 1.71 1.75 3.045 ;
        RECT 1.49 0.395 1.75 1.04 ;
        RECT 0.635 1.71 0.89 3.045 ;
        RECT 0.175 0.84 0.345 1.885 ;
    END
  END Y
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.69 5.69 2.945 ;
      LAYER li ;
        RECT 5.36 2.055 5.615 3.075 ;
        RECT 4.5 2.055 4.76 3.075 ;
        RECT 3.64 2.055 3.9 3.075 ;
        RECT 2.78 2.055 3.04 3.075 ;
        RECT 1.92 2.055 2.18 3.075 ;
        RECT 1.06 2.055 1.32 3.075 ;
        RECT 0.2 2.055 0.46 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.5 -0.085 4.795 0.67 ;
        RECT 3.64 -0.085 3.9 0.67 ;
        RECT 2.78 -0.085 3.04 0.67 ;
        RECT 1.92 -0.085 2.18 0.67 ;
        RECT 1.025 -0.085 1.32 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_invkapwr_8

MACRO scs130lp_invlp_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invlp_0 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 2.15 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3021 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 2.32 1.315 3 ;
        RECT 1.085 0.44 1.315 3 ;
        RECT 0.985 0.44 1.315 0.9 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.165 -0.085 0.495 0.9 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.165 2.32 0.495 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_invlp_0

MACRO scs130lp_invlp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invlp_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.455 1.515 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.255 1.315 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.165 -0.085 0.495 1.01 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.195 1.815 0.525 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_invlp_1

MACRO scs130lp_invlp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invlp_2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.455 1.555 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.595 1.315 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.995 -0.085 2.245 1.135 ;
        RECT 0.125 -0.085 0.455 1.01 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.915 1.815 2.245 3.415 ;
        RECT 0.125 1.815 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.485 0.255 1.815 1.135 ;
      RECT 0.635 0.255 0.805 1.135 ;
      RECT 0.635 0.255 1.815 0.425 ;
      RECT 0.635 2.905 1.745 3.075 ;
      RECT 1.495 1.815 1.745 3.075 ;
      RECT 0.635 1.815 0.805 3.075 ;
  END
END scs130lp_invlp_2

MACRO scs130lp_invlp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invlp_4 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.385 1.345 4.095 1.675 ;
        RECT 1.565 1.345 2.755 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4112 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.925 1.845 3.255 2.735 ;
        RECT 1.045 1.005 3.235 1.175 ;
        RECT 2.905 0.595 3.235 1.175 ;
        RECT 1.045 1.95 3.255 2.12 ;
        RECT 1.925 1.95 2.255 2.735 ;
        RECT 2.055 0.595 2.225 1.175 ;
        RECT 1.045 1.005 1.215 2.12 ;
        RECT 0.605 1.18 1.215 1.41 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.915 -0.085 4.165 1.125 ;
        RECT 1.045 -0.085 1.375 0.495 ;
        RECT 0.115 -0.085 0.365 1.125 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.855 1.845 4.185 3.415 ;
        RECT 0.995 2.63 1.245 3.415 ;
        RECT 0.135 1.815 0.385 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.405 0.255 3.735 1.125 ;
      RECT 0.545 0.255 0.875 1.01 ;
      RECT 2.405 0.255 2.735 0.835 ;
      RECT 0.545 0.665 1.875 0.835 ;
      RECT 1.545 0.255 1.875 0.835 ;
      RECT 1.545 0.255 3.735 0.425 ;
      RECT 1.425 2.905 3.685 3.075 ;
      RECT 3.435 1.845 3.685 3.075 ;
      RECT 0.565 1.815 0.815 3.075 ;
      RECT 2.425 2.29 2.755 3.075 ;
      RECT 1.425 2.29 1.755 3.075 ;
      RECT 0.565 2.29 1.755 2.46 ;
  END
END scs130lp_invlp_4

MACRO scs130lp_invlp_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invlp_8 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 5.04 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.305 1.345 7.415 1.675 ;
        RECT 1.565 1.345 3.235 1.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.499 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.345 1.845 6.675 2.735 ;
        RECT 0.965 1.005 6.605 1.175 ;
        RECT 6.275 0.595 6.605 1.175 ;
        RECT 3.775 1.845 6.675 2.015 ;
        RECT 5.495 1.845 5.665 2.735 ;
        RECT 5.275 0.595 5.605 1.175 ;
        RECT 4.635 1.845 4.805 2.735 ;
        RECT 4.495 0.595 4.745 1.175 ;
        RECT 3.775 1.845 3.945 2.735 ;
        RECT 3.555 0.595 3.805 1.175 ;
        RECT 0.965 1.95 3.945 2.12 ;
        RECT 0.965 1.005 1.135 2.12 ;
        RECT 0.605 1.55 1.135 1.78 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.285 -0.085 7.535 1.125 ;
        RECT 2.695 -0.085 3.025 0.495 ;
        RECT 1.835 -0.085 2.165 0.495 ;
        RECT 0.975 -0.085 1.305 0.495 ;
        RECT 0.115 -0.085 0.365 1.125 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.205 1.845 7.535 3.415 ;
        RECT 2.765 2.63 3.095 3.415 ;
        RECT 1.835 2.63 2.085 3.415 ;
        RECT 0.975 2.63 1.305 3.415 ;
        RECT 0.115 1.815 0.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.775 0.255 7.105 1.125 ;
      RECT 0.545 0.255 0.795 1.125 ;
      RECT 5.775 0.255 6.105 0.835 ;
      RECT 4.925 0.255 5.095 0.835 ;
      RECT 3.985 0.255 4.315 0.835 ;
      RECT 0.545 0.665 3.375 0.835 ;
      RECT 3.205 0.255 3.375 0.835 ;
      RECT 2.345 0.255 2.515 0.835 ;
      RECT 1.485 0.255 1.655 0.835 ;
      RECT 3.205 0.255 7.105 0.425 ;
      RECT 3.265 2.905 7.025 3.075 ;
      RECT 6.855 1.845 7.025 3.075 ;
      RECT 2.265 2.29 2.595 3.075 ;
      RECT 1.485 2.29 1.655 3.075 ;
      RECT 0.545 1.95 0.795 3.075 ;
      RECT 5.845 2.185 6.175 3.075 ;
      RECT 4.985 2.185 5.315 3.075 ;
      RECT 4.125 2.185 4.455 3.075 ;
      RECT 3.265 2.29 3.595 3.075 ;
      RECT 0.545 2.29 3.595 2.46 ;
  END
END scs130lp_invlp_8

MACRO scs130lp_invlp_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_invlp_m 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 2.15 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 2.43 1.315 2.89 ;
        RECT 1.085 0.44 1.315 2.89 ;
        RECT 0.985 0.44 1.315 0.9 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.165 -0.085 0.495 0.9 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.165 2.43 0.495 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_invlp_m

MACRO scs130lp_iso0n_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso0n_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.345 1.395 1.09 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.855 0.465 3.275 3.075 ;
    END
  END X
  PIN sleepb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.315 1.395 1.985 1.75 ;
    END
  END sleepb
  PIN kagnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.07 0.44 3.29 0.67 ;
      LAYER li ;
        RECT 1.44 0.39 2.275 0.84 ;
    END
  END kagnd
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.99 2.295 2.675 3.415 ;
        RECT 0.29 2.49 0.62 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.08 1.955 1.41 2.82 ;
      RECT 1.08 1.955 2.685 2.125 ;
      RECT 2.275 1.055 2.685 2.125 ;
      RECT 0.65 1.055 2.685 1.225 ;
      RECT 0.65 0.51 0.98 1.225 ;
  END
END scs130lp_iso0n_lp

MACRO scs130lp_iso0n_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso0n_lp2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.955 0.455 1.78 ;
    END
  END A
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 1.515 1.795 1.845 ;
    END
  END SLEEPB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.795 2.025 2.275 3.065 ;
        RECT 2.045 0.305 2.275 3.065 ;
        RECT 1.945 0.305 2.275 0.765 ;
    END
  END X
  PIN kagnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.07 0.44 2.33 0.67 ;
      LAYER li ;
        RECT 1.085 0.305 1.455 0.765 ;
    END
  END kagnd
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.265 2.025 1.595 3.415 ;
        RECT 0.14 2.025 0.47 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.65 2.025 1.065 3.065 ;
      RECT 0.65 0.595 0.82 3.065 ;
      RECT 0.65 0.945 1.72 1.275 ;
      RECT 0.305 0.595 0.82 0.765 ;
      RECT 0.305 0.305 0.635 0.765 ;
  END
END scs130lp_iso0n_lp2

MACRO scs130lp_iso0p_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso0p_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 1.395 2.65 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.4 0.465 3.755 3.075 ;
    END
  END X
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 1.16 0.92 1.895 ;
    END
  END sleep
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.66 3.77 2.89 ;
      LAYER li ;
        RECT 2.525 2.295 2.91 3.075 ;
        RECT 0.895 2.445 1.225 2.92 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.55 -0.085 2.885 0.835 ;
        RECT 0.895 -0.085 1.575 0.84 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.765 1.955 1.975 2.855 ;
      RECT 1.765 1.955 3.23 2.125 ;
      RECT 2.82 1.005 3.23 2.125 ;
      RECT 2.095 1.005 3.23 1.225 ;
      RECT 2.095 0.43 2.305 1.225 ;
      RECT 0.155 0.43 0.375 2.855 ;
      RECT 0.155 2.065 1.595 2.235 ;
      RECT 1.2 1.39 1.595 2.235 ;
  END
END scs130lp_iso0p_lp

MACRO scs130lp_iso0p_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso0p_lp2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 1.395 2.755 1.75 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 1.01 0.92 1.78 ;
    END
  END SLEEP
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3763 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.4 0.465 3.755 3.075 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.66 3.77 2.89 ;
      LAYER li ;
        RECT 2.235 2.295 3.145 3.075 ;
        RECT 0.635 2.29 1.485 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.55 -0.085 2.885 0.835 ;
        RECT 0.895 -0.085 1.575 0.84 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.765 1.955 1.975 3.075 ;
      RECT 1.765 1.955 3.23 2.125 ;
      RECT 2.925 1.005 3.23 2.125 ;
      RECT 2.095 1.005 3.23 1.225 ;
      RECT 2.095 0.43 2.305 1.225 ;
      RECT 0.155 0.43 0.375 3.075 ;
      RECT 0.155 1.95 1.595 2.12 ;
      RECT 1.2 1.01 1.595 2.12 ;
  END
END scs130lp_iso0p_lp2

MACRO scs130lp_iso1n_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso1n_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.91 1.395 2.58 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.395 0.465 3.755 3.075 ;
    END
  END X
  PIN sleepb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.54 1.16 1.16 1.99 ;
    END
  END sleepb
  PIN kagnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.07 0.44 3.77 0.67 ;
      LAYER li ;
        RECT 2.525 0.43 3.155 0.885 ;
        RECT 0.885 0.43 1.515 0.885 ;
    END
  END kagnd
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.525 2.295 2.91 3.415 ;
        RECT 1.19 2.5 1.52 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.095 1.955 2.305 2.88 ;
      RECT 2.095 1.955 3.225 2.125 ;
      RECT 2.895 1.055 3.225 2.125 ;
      RECT 1.87 1.055 3.225 1.225 ;
      RECT 1.87 0.43 2.065 1.225 ;
      RECT 1.735 0.43 2.065 0.885 ;
      RECT 0.345 2.16 0.59 2.82 ;
      RECT 0.125 2.16 1.7 2.33 ;
      RECT 1.37 1.315 1.7 2.33 ;
      RECT 0.125 0.885 0.37 2.33 ;
      RECT 0.12 0.43 0.365 0.885 ;
  END
END scs130lp_iso1n_lp

MACRO scs130lp_iso1n_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso1n_lp2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.165 2.755 1.495 ;
    END
  END A
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.505 1.515 0.835 1.845 ;
    END
  END SLEEPB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 2.025 3.715 3.065 ;
        RECT 3.435 0.525 3.715 3.065 ;
        RECT 3.385 0.525 3.715 0.985 ;
    END
  END X
  PIN kagnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.07 0.44 3.77 0.67 ;
      LAYER li ;
        RECT 2.445 0.265 3.075 0.985 ;
        RECT 0.755 0.265 3.075 0.435 ;
        RECT 0.755 0.265 1.385 0.985 ;
    END
  END kagnd
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.855 2.025 3.185 3.415 ;
        RECT 0.905 2.025 1.235 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.695 1.675 2.295 3.065 ;
      RECT 1.695 1.675 3.265 1.845 ;
      RECT 2.935 1.175 3.265 1.845 ;
      RECT 1.695 0.615 1.865 3.065 ;
      RECT 1.695 0.615 2.055 0.985 ;
      RECT 0.115 2.025 0.625 3.065 ;
      RECT 0.115 0.525 0.285 3.065 ;
      RECT 1.17 1.165 1.5 1.835 ;
      RECT 0.115 1.165 1.5 1.335 ;
      RECT 0.115 0.525 0.445 1.335 ;
  END
END scs130lp_iso1n_lp2

MACRO scs130lp_iso1p_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso1p_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 1.35 1.225 1.75 ;
        RECT 0.555 1.16 0.855 1.75 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4452 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.855 0.465 3.275 3.075 ;
    END
  END X
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.435 1.35 2.105 1.75 ;
    END
  END sleep
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.66 3.29 2.89 ;
      LAYER li ;
        RECT 1.56 2.295 2.365 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.01 -0.085 2.34 0.84 ;
        RECT 0.46 -0.085 0.76 0.84 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.77 1.955 1.1 2.82 ;
      RECT 0.77 1.955 2.685 2.125 ;
      RECT 2.35 1.01 2.685 2.125 ;
      RECT 1.28 1.01 2.685 1.18 ;
      RECT 1.28 0.44 1.49 1.18 ;
  END
END scs130lp_iso1p_lp

MACRO scs130lp_iso1p_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_iso1p_lp2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.005 0.915 1.78 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.16 1.795 1.83 ;
    END
  END SLEEP
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.71 0.265 3.235 2.52 ;
        RECT 2.505 1.92 2.835 3.065 ;
    END
  END X
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.66 3.29 2.89 ;
      LAYER li ;
        RECT 1.635 2.025 2.335 3.065 ;
        RECT 1.345 2.66 2.335 2.89 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.89 -0.085 2.22 0.64 ;
        RECT 0.28 -0.085 0.61 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.645 2.025 0.975 3.065 ;
      RECT 0.645 2.025 1.27 2.195 ;
      RECT 1.1 0.265 1.27 2.195 ;
      RECT 2.195 0.82 2.525 1.535 ;
      RECT 1.1 0.82 2.525 0.99 ;
      RECT 1.1 0.265 1.43 0.99 ;
  END
END scs130lp_iso1p_lp2

MACRO scs130lp_isobufsrc_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_isobufsrc_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.425 0.865 1.75 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.425 1.415 1.75 ;
    END
  END SLEEP
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8526 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.925 1.815 2.315 3.075 ;
        RECT 2.055 0.745 2.315 3.075 ;
        RECT 1.39 0.745 2.315 0.915 ;
        RECT 1.39 0.255 1.65 0.915 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.82 -0.085 2.15 0.575 ;
        RECT 0.795 -0.085 1.22 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.96 2.31 1.29 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.42 1.92 1.755 2.14 ;
      RECT 1.585 1.085 1.755 2.14 ;
      RECT 1.585 1.085 1.885 1.515 ;
      RECT 0.355 1.085 1.885 1.255 ;
      RECT 0.355 0.285 0.625 1.255 ;
  END
END scs130lp_isobufsrc_1

MACRO scs130lp_isobufsrc_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_isobufsrc_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 1.185 0.885 1.515 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.075 2.815 1.515 ;
        RECT 1.055 1.075 2.815 1.245 ;
        RECT 1.055 1.075 1.775 1.435 ;
    END
  END SLEEP
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8232 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.82 2.025 3.275 2.195 ;
        RECT 2.985 0.735 3.275 2.195 ;
        RECT 1.435 0.735 3.275 0.905 ;
        RECT 2.365 0.255 2.555 0.905 ;
        RECT 1.82 2.025 2.15 2.715 ;
        RECT 1.435 0.255 1.695 0.905 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.725 -0.085 3.055 0.565 ;
        RECT 1.865 -0.085 2.195 0.565 ;
        RECT 0.62 -0.085 1.265 0.885 ;
        RECT 0.62 -0.085 0.895 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.68 2.365 3.01 3.415 ;
        RECT 0.865 2.025 1.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.42 2.895 2.51 3.075 ;
      RECT 2.32 2.365 2.51 3.075 ;
      RECT 1.42 2.025 1.65 3.075 ;
      RECT 0.16 1.685 0.695 2.21 ;
      RECT 0.16 1.685 2.275 1.855 ;
      RECT 1.945 1.415 2.275 1.855 ;
      RECT 0.16 0.7 0.43 2.21 ;
  END
END scs130lp_isobufsrc_2

MACRO scs130lp_isobufsrc_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_isobufsrc_4 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.345 0.435 1.76 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.965 1.695 4.305 1.865 ;
        RECT 4.045 1.345 4.305 1.865 ;
        RECT 2.065 1.425 3.205 1.865 ;
        RECT 0.965 1.425 1.295 1.865 ;
    END
  END SLEEP
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.63 2.035 4.7 2.205 ;
        RECT 4.475 1.005 4.7 2.205 ;
        RECT 3.84 1.005 4.7 1.175 ;
        RECT 3.84 0.745 4.03 1.175 ;
        RECT 3.85 0.255 4.03 1.175 ;
        RECT 1.2 0.745 4.03 0.915 ;
        RECT 3.41 2.035 3.62 2.715 ;
        RECT 2.92 0.255 3.25 0.915 ;
        RECT 2.06 0.255 2.39 0.915 ;
        RECT 1.63 2.035 1.96 2.255 ;
        RECT 1.2 0.255 1.53 0.915 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.21 -0.085 4.54 0.835 ;
        RECT 3.42 -0.085 3.68 0.575 ;
        RECT 2.56 -0.085 2.75 0.575 ;
        RECT 1.7 -0.085 1.89 0.575 ;
        RECT 0.69 -0.085 1.02 0.835 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.21 2.375 4.54 3.415 ;
        RECT 0.75 2.425 2.82 2.655 ;
        RECT 0.75 2.27 1.08 2.655 ;
        RECT 0.75 2.27 1.03 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.2 2.885 4.04 3.065 ;
      RECT 3.84 2.375 4.04 3.065 ;
      RECT 1.2 2.825 3.19 3.065 ;
      RECT 2.99 2.375 3.19 3.065 ;
      RECT 0.26 1.93 0.53 3.075 ;
      RECT 0.26 1.93 0.785 2.1 ;
      RECT 0.615 1.005 0.785 2.1 ;
      RECT 3.375 1.085 3.635 1.515 ;
      RECT 1.565 1.085 1.895 1.515 ;
      RECT 0.615 1.085 3.635 1.255 ;
      RECT 0.26 1.005 0.785 1.175 ;
      RECT 0.26 0.255 0.52 1.175 ;
  END
END scs130lp_isobufsrc_4

MACRO scs130lp_isolatch_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_isolatch_lp 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.255 0.835 1.78 ;
        RECT 0.125 2.185 0.585 2.515 ;
        RECT 0.125 1.255 0.295 2.515 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4597 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.45 0.44 7.085 2.955 ;
    END
  END Q
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.355 1.45 4.685 1.78 ;
    END
  END SLEEPB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 7.13 2.945 ;
      LAYER li ;
        RECT 5.865 1.915 6.195 2.955 ;
        RECT 4.775 2.29 5.155 2.905 ;
        RECT 2.515 2.125 2.845 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 5.95 -0.085 6.28 1.325 ;
        RECT 4.6 -0.085 4.85 0.905 ;
        RECT 2.97 -0.085 3.22 0.775 ;
        RECT 0.59 -0.085 0.92 0.745 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 0.13 2.685 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.515 2.905 4.605 3.075 ;
      RECT 4.435 1.95 4.605 3.075 ;
      RECT 5.335 1.915 5.665 2.955 ;
      RECT 5.495 0.445 5.665 2.955 ;
      RECT 3.515 1.785 3.845 3.075 ;
      RECT 4.435 1.95 5.665 2.12 ;
      RECT 5.46 0.445 5.665 0.775 ;
      RECT 1.495 2.29 1.855 2.735 ;
      RECT 1.685 1.33 1.855 2.735 ;
      RECT 4.895 1.075 5.225 1.745 ;
      RECT 1.575 0.345 1.745 1.5 ;
      RECT 4.15 1.075 5.225 1.245 ;
      RECT 2.415 0.945 3.56 1.115 ;
      RECT 3.39 0.255 3.56 1.115 ;
      RECT 4.15 0.255 4.32 1.245 ;
      RECT 2.415 0.555 2.585 1.115 ;
      RECT 1.575 0.555 2.585 0.725 ;
      RECT 1.575 0.345 1.97 0.725 ;
      RECT 3.39 0.255 4.32 0.425 ;
      RECT 4.015 2.055 4.265 2.735 ;
      RECT 4.015 1.445 4.185 2.735 ;
      RECT 2.075 1.445 4.185 1.615 ;
      RECT 2.075 1.285 3.98 1.615 ;
      RECT 3.73 0.595 3.98 1.615 ;
      RECT 2.075 0.895 2.245 1.615 ;
      RECT 1.915 0.895 2.245 1.16 ;
      RECT 3.045 1.785 3.295 3.075 ;
      RECT 1.155 2.905 2.345 3.075 ;
      RECT 2.175 1.785 2.345 3.075 ;
      RECT 1.155 1.95 1.325 3.075 ;
      RECT 1.185 1.67 1.515 2.12 ;
      RECT 2.175 1.785 3.295 1.955 ;
      RECT 1.185 0.915 1.355 2.12 ;
      RECT 0.16 0.915 1.355 1.085 ;
      RECT 0.16 0.345 0.41 1.085 ;
  END
END scs130lp_isolatch_lp

MACRO scs130lp_lsbuf_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_lsbuf_lp 0 0 ;
  SIZE 4.8 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.678 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.075 2.775 1.91 3.075 ;
        RECT 1.075 1.53 1.245 3.075 ;
        RECT 0.585 1.53 1.245 2.135 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4876 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.895 3.585 4.225 6.405 ;
    END
  END X
  PIN destvpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 5.22 0.39 6.395 ;
    END
    PORT
      LAYER li ;
        RECT 4.41 5.22 4.71 6.395 ;
    END
  END destvpb
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 0.265 0.39 1.44 ;
    END
    PORT
      LAYER li ;
        RECT 4.41 0.265 4.71 1.44 ;
    END
  END vpb
  PIN destpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 6.415 4.8 6.905 ;
      LAYER li ;
        RECT 0 6.575 4.8 6.745 ;
        RECT 3.105 5.5 3.435 6.745 ;
        RECT 1.715 5.695 2.045 6.745 ;
    END
  END destpwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 2.505 3.245 4.8 3.415 ;
        RECT 4.41 1.89 4.71 4.77 ;
        RECT 3.105 3.245 3.435 4.23 ;
        RECT 1.715 3.245 1.995 4.48 ;
        RECT 0 3.245 1.995 3.415 ;
        RECT 0.575 2.305 0.905 3.415 ;
        RECT 0.09 1.89 0.39 4.77 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 0.575 -0.085 0.905 1.175 ;
    END
  END vpwr
  OBS
    LAYER li ;
      RECT 2.505 5.355 2.835 6.395 ;
      RECT 2.665 5.16 2.835 6.395 ;
      RECT 1.51 5.355 2.835 5.525 ;
      RECT 1.51 4.99 1.68 5.525 ;
      RECT 2.665 5.16 3.16 5.33 ;
      RECT 2.99 4.4 3.16 5.33 ;
      RECT 1.35 4.99 1.68 5.265 ;
      RECT 2.765 4.4 3.16 4.57 ;
      RECT 2.55 3.585 2.935 4.44 ;
      RECT 2.505 3.585 2.935 4.14 ;
      RECT 2.45 4.74 2.82 4.99 ;
      RECT 2.21 4.61 2.595 4.84 ;
      RECT 2.21 4.31 2.38 4.84 ;
      RECT 2.165 2.435 2.335 4.48 ;
      RECT 1.415 2.435 2.335 2.605 ;
      RECT 1.415 0.265 1.715 2.605 ;
      RECT 1.365 0.265 1.715 1.36 ;
      RECT 0.925 5.435 1.275 6.405 ;
      RECT 0.925 3.585 1.18 6.405 ;
      RECT 1.87 5.01 2.28 5.185 ;
      RECT 1.87 4.65 2.04 5.185 ;
      RECT 0.925 4.65 2.04 4.82 ;
      RECT 0.925 3.585 1.205 4.82 ;
  END
END scs130lp_lsbuf_lp

MACRO scs130lp_lsbufiso0p_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_lsbufiso0p_lp 0 0 ;
  SIZE 6.72 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.678 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.075 2.775 1.645 3.075 ;
        RECT 1.075 1.53 1.245 3.075 ;
        RECT 0.585 1.53 1.245 2.135 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7144 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.815 3.585 6.145 6.405 ;
        RECT 4.285 4.32 6.145 4.49 ;
        RECT 4.285 3.59 4.565 4.49 ;
    END
  END X
  PIN destvpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 5.22 0.39 6.395 ;
    END
    PORT
      LAYER li ;
        RECT 6.33 5.22 6.63 6.395 ;
    END
  END destvpb
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.978 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.835 4.505 3.42 4.91 ;
    END
  END sleep
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 0.265 0.39 1.44 ;
    END
    PORT
      LAYER li ;
        RECT 6.33 0.265 6.63 1.44 ;
    END
  END vpb
  PIN destpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 6.415 6.72 6.905 ;
      LAYER li ;
        RECT 0 6.575 6.72 6.745 ;
        RECT 5.04 5.42 5.355 6.745 ;
        RECT 3.57 5.42 3.74 6.745 ;
    END
  END destpwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 3.075 6.72 3.565 ;
      LAYER li ;
        RECT 2.7 3.245 6.72 3.415 ;
        RECT 6.33 1.89 6.63 4.77 ;
        RECT 5.025 3.245 5.355 3.88 ;
        RECT 2.71 2.43 3.04 3.415 ;
        RECT 2.7 3.245 3.03 4.24 ;
        RECT 0 3.245 2.145 3.415 ;
        RECT 0.575 2.305 0.905 3.415 ;
        RECT 0.09 1.89 0.39 4.77 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 0.575 -0.085 0.905 1.175 ;
    END
  END vpwr
  OBS
    LAYER li ;
      RECT 3.99 6.235 4.87 6.405 ;
      RECT 4.7 4.66 4.87 6.405 ;
      RECT 3.99 5.08 4.16 6.405 ;
      RECT 2.495 5.08 2.745 5.295 ;
      RECT 2.495 5.08 4.16 5.25 ;
      RECT 2.495 4.935 2.665 5.295 ;
      RECT 4.7 4.66 5.58 4.99 ;
      RECT 4.33 4.74 4.53 6.055 ;
      RECT 3.59 4.74 4.53 4.91 ;
      RECT 3.59 3.585 3.815 4.91 ;
      RECT 3.49 3.585 3.82 4.24 ;
      RECT 3.49 3.585 4.08 3.915 ;
      RECT 1.365 6.235 3.39 6.405 ;
      RECT 3.06 5.465 3.39 6.405 ;
      RECT 1.365 5.695 1.695 6.405 ;
      RECT 1.365 3.585 1.645 4.48 ;
      RECT 1.365 3.585 2.485 3.755 ;
      RECT 2.315 2.33 2.485 3.755 ;
      RECT 2.315 2.33 2.53 3.09 ;
      RECT 2.155 5.465 2.485 6.055 ;
      RECT 1.16 5.355 2.325 5.525 ;
      RECT 2.155 4.07 2.325 6.055 ;
      RECT 1.16 4.99 1.33 5.525 ;
      RECT 1 4.99 1.33 5.265 ;
      RECT 2.155 4.07 2.485 4.4 ;
      RECT 1.815 2.435 2.145 3.075 ;
      RECT 1.415 2.435 2.145 2.605 ;
      RECT 1.415 0.265 1.715 2.605 ;
      RECT 1.365 0.265 1.715 1.36 ;
      RECT 0.575 5.435 0.925 6.405 ;
      RECT 0.575 3.585 0.83 6.405 ;
      RECT 1.52 5.01 1.93 5.185 ;
      RECT 1.52 4.65 1.69 5.185 ;
      RECT 0.575 4.65 1.69 4.82 ;
      RECT 0.575 3.585 0.855 4.82 ;
  END
END scs130lp_lsbufiso0p_lp

MACRO scs130lp_lsbufiso1p_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_lsbufiso1p_lp 0 0 ;
  SIZE 7.2 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.678 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.075 2.775 1.645 3.075 ;
        RECT 1.075 1.53 1.245 3.075 ;
        RECT 0.585 1.53 1.245 2.135 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7726 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.29 3.585 6.62 6.405 ;
        RECT 4.71 5.42 6.62 5.59 ;
        RECT 4.71 5.42 5.04 6.405 ;
    END
  END X
  PIN destvpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 5.22 0.39 6.395 ;
    END
    PORT
      LAYER li ;
        RECT 6.81 5.22 7.11 6.395 ;
    END
  END destvpb
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.576 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.835 4.505 3.42 4.91 ;
    END
  END sleep
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 0.265 0.39 1.44 ;
    END
    PORT
      LAYER li ;
        RECT 6.81 0.265 7.11 1.44 ;
    END
  END vpb
  PIN destpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 6.415 7.2 6.905 ;
      LAYER li ;
        RECT 0 6.575 7.2 6.745 ;
        RECT 5.5 5.76 5.83 6.745 ;
        RECT 3.21 5.455 3.38 6.745 ;
    END
  END destpwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 3.075 7.2 3.565 ;
      LAYER li ;
        RECT 2.7 3.245 7.2 3.415 ;
        RECT 6.81 1.89 7.11 4.77 ;
        RECT 5.5 3.245 5.83 4.23 ;
        RECT 2.7 2.43 3.04 3.415 ;
        RECT 2.7 2.43 3.03 4.24 ;
        RECT 0 3.245 2.145 3.415 ;
        RECT 0.575 2.305 0.905 3.415 ;
        RECT 0.09 1.89 0.39 4.77 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 0.575 -0.085 0.905 1.175 ;
    END
  END vpwr
  OBS
    LAYER li ;
      RECT 3.63 6.235 4.515 6.405 ;
      RECT 4.34 4.865 4.515 6.405 ;
      RECT 3.63 5.08 3.8 6.405 ;
      RECT 2.495 5.08 3.8 5.285 ;
      RECT 4.34 4.865 6.055 5.195 ;
      RECT 2.495 4.935 2.665 5.285 ;
      RECT 3.97 4.74 4.17 6.055 ;
      RECT 3.59 4.74 4.17 4.91 ;
      RECT 3.59 3.585 3.815 4.91 ;
      RECT 3.49 3.585 3.82 4.24 ;
      RECT 3.49 3.585 4.08 3.915 ;
      RECT 1.365 6.235 3.03 6.405 ;
      RECT 2.7 5.465 3.03 6.405 ;
      RECT 1.365 5.695 1.695 6.405 ;
      RECT 1.365 3.585 1.645 4.48 ;
      RECT 1.365 3.585 2.485 3.755 ;
      RECT 2.315 2.33 2.485 3.755 ;
      RECT 2.315 2.33 2.53 3.09 ;
      RECT 2.155 5.465 2.485 6.055 ;
      RECT 1.16 5.355 2.325 5.525 ;
      RECT 2.155 4.07 2.325 6.055 ;
      RECT 1.16 4.99 1.33 5.525 ;
      RECT 1 4.99 1.33 5.265 ;
      RECT 2.155 4.07 2.485 4.4 ;
      RECT 1.815 2.435 2.145 3.075 ;
      RECT 1.415 2.435 2.145 2.605 ;
      RECT 1.415 0.265 1.715 2.605 ;
      RECT 1.365 0.265 1.715 1.36 ;
      RECT 0.575 5.435 0.925 6.405 ;
      RECT 0.575 3.585 0.83 6.405 ;
      RECT 1.52 5.01 1.93 5.185 ;
      RECT 1.52 4.65 1.69 5.185 ;
      RECT 0.575 4.65 1.69 4.82 ;
      RECT 0.575 3.585 0.855 4.82 ;
  END
END scs130lp_lsbufiso1p_lp

MACRO scs130lp_maj3_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_maj3_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 0.905 1.515 1.575 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 0.905 2.755 1.575 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 2.66 2.925 3.065 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3757 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.465 0.265 3.715 2.595 ;
        RECT 3.15 0.265 3.715 0.725 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.72 -0.085 2.97 0.725 ;
        RECT 1.11 -0.085 1.44 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.105 2.105 3.275 3.415 ;
        RECT 2.84 2.105 3.275 2.48 ;
        RECT 1.025 2.135 1.355 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.93 1.755 2.26 2.595 ;
      RECT 0.12 1.755 0.45 2.595 ;
      RECT 0.12 1.755 3.285 1.925 ;
      RECT 2.955 1.105 3.285 1.925 ;
      RECT 1.695 0.265 1.865 1.925 ;
      RECT 0.12 0.265 0.29 2.595 ;
      RECT 1.695 0.265 2.26 0.725 ;
      RECT 0.12 0.265 0.62 0.725 ;
  END
END scs130lp_maj3_0

MACRO scs130lp_maj3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_maj3_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.125 1.375 1.455 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.18 2.275 1.51 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 2.66 2.755 3.065 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.475 0.265 3.725 3.065 ;
        RECT 3.355 0.265 3.725 1.145 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.845 -0.085 3.175 1.145 ;
        RECT 1.07 -0.085 1.4 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.965 1.835 3.295 3.415 ;
        RECT 0.92 1.935 1.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.825 1.925 2.155 2.395 ;
      RECT 0.13 1.935 0.46 2.395 ;
      RECT 1.825 1.925 2.625 2.095 ;
      RECT 2.455 0.265 2.625 2.095 ;
      RECT 0.13 0.265 0.3 2.395 ;
      RECT 2.455 1.325 3.295 1.655 ;
      RECT 0.13 0.775 2.625 0.945 ;
      RECT 1.94 0.265 2.625 0.945 ;
      RECT 0.13 0.265 0.38 0.945 ;
      RECT 0.56 0.265 0.89 0.595 ;
  END
END scs130lp_maj3_1

MACRO scs130lp_maj3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_maj3_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.215 1.795 1.885 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 1.215 2.31 1.885 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 2.065 3.235 2.235 ;
        RECT 2.525 1.905 3.235 2.235 ;
        RECT 0.44 1.265 0.77 2.235 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.445 1.795 3.775 3.065 ;
        RECT 3.605 0.265 3.775 3.065 ;
        RECT 3.285 0.265 3.775 1.105 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.955 -0.085 4.205 1.105 ;
        RECT 2.775 -0.085 3.105 0.685 ;
        RECT 1.135 -0.085 1.465 0.685 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.955 1.795 4.205 3.415 ;
        RECT 2.735 2.415 3.065 3.415 ;
        RECT 1.095 2.765 1.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.915 2.415 2.245 3.065 ;
      RECT 0.09 2.415 0.605 3.065 ;
      RECT 0.09 2.415 2.245 2.585 ;
      RECT 0.09 0.865 0.26 3.065 ;
      RECT 2.935 1.285 3.425 1.615 ;
      RECT 2.935 0.865 3.105 1.615 ;
      RECT 0.09 0.865 3.105 1.035 ;
      RECT 1.955 0.265 2.285 1.035 ;
      RECT 0.315 0.265 0.645 1.035 ;
  END
END scs130lp_maj3_2

MACRO scs130lp_maj3_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_maj3_4 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.18 1.415 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.18 2.305 1.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.485 1.275 2.98 1.605 ;
        RECT 0.735 2.225 2.655 2.395 ;
        RECT 2.485 1.275 2.655 2.395 ;
        RECT 0.735 1.18 0.905 2.395 ;
        RECT 0.44 1.18 0.905 1.515 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2096 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.345 1.785 5.155 1.955 ;
        RECT 4.925 0.925 5.155 1.955 ;
        RECT 3.51 0.925 5.155 1.095 ;
        RECT 4.365 1.785 4.695 3.065 ;
        RECT 4.325 0.265 4.655 1.095 ;
        RECT 3.51 0.265 3.68 1.095 ;
        RECT 3.345 1.785 3.675 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.835 -0.085 5.165 0.745 ;
        RECT 3.86 -0.085 4.11 0.745 ;
        RECT 2.775 -0.085 3.105 0.65 ;
        RECT 1.135 -0.085 1.465 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.875 2.135 5.125 3.415 ;
        RECT 3.855 2.135 4.185 3.415 ;
        RECT 2.835 1.795 3.165 3.415 ;
        RECT 1.135 2.575 1.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.09 1.795 0.555 3.065 ;
      RECT 1.625 1.795 2.285 2.045 ;
      RECT 1.625 0.83 1.795 2.045 ;
      RECT 0.09 0.83 0.26 3.065 ;
      RECT 3.16 1.275 4.67 1.605 ;
      RECT 3.16 0.83 3.33 1.605 ;
      RECT 0.09 0.83 3.33 1 ;
      RECT 1.955 0.295 2.285 1 ;
      RECT 0.315 0.265 0.645 1 ;
  END
END scs130lp_maj3_4

MACRO scs130lp_maj3_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_maj3_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.605 1.795 2.15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.42 1.245 2.75 1.915 ;
        RECT 0.44 1.245 2.75 1.415 ;
        RECT 0.44 1.225 1.315 1.415 ;
        RECT 1.085 1.18 1.315 1.415 ;
        RECT 0.44 1.225 0.76 1.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.96 1.245 3.29 1.915 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.755 1.92 4.21 3.065 ;
        RECT 4.04 0.32 4.21 3.065 ;
        RECT 3.875 0.32 4.21 0.78 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.085 -0.085 3.415 0.715 ;
        RECT 1.215 -0.085 1.545 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.215 2.095 3.545 3.415 ;
        RECT 1.195 2.68 1.525 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.185 2.095 2.515 3.065 ;
      RECT 0.09 2.075 0.455 3.065 ;
      RECT 0.09 2.33 2.515 2.5 ;
      RECT 0.09 0.875 0.26 3.065 ;
      RECT 3.525 0.985 3.86 1.655 ;
      RECT 1.495 0.895 3.695 1.065 ;
      RECT 0.09 0.875 0.645 1.045 ;
      RECT 0.315 0.605 0.645 1.045 ;
      RECT 0.315 0.83 1.665 1 ;
      RECT 2.195 0.32 2.525 1.065 ;
  END
END scs130lp_maj3_lp

MACRO scs130lp_maj3_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_maj3_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 0.905 1.325 1.575 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.905 2.275 1.575 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.455 2.29 2.785 3.065 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.395 0.265 3.725 2.89 ;
        RECT 3.315 0.265 3.725 0.725 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.805 -0.085 3.135 0.725 ;
        RECT 0.97 -0.085 1.3 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.965 2.105 3.215 3.415 ;
        RECT 0.97 2.105 1.3 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.79 1.755 2.12 2.565 ;
      RECT 0.15 1.755 0.48 2.565 ;
      RECT 0.15 1.755 3.215 1.925 ;
      RECT 2.885 1.255 3.215 1.925 ;
      RECT 2.455 0.555 2.625 1.925 ;
      RECT 0.15 0.265 0.32 2.565 ;
      RECT 1.79 0.555 2.625 0.725 ;
      RECT 0.15 0.265 0.48 0.725 ;
      RECT 1.79 0.265 2.12 0.725 ;
  END
END scs130lp_maj3_m

MACRO scs130lp_mux2_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 1.21 1.775 1.645 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 2.155 2.465 2.705 ;
        RECT 2.295 0.265 2.465 2.705 ;
        RECT 1.645 0.265 2.465 0.5 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.635 2.32 3.385 2.49 ;
        RECT 2.985 1.515 3.385 2.49 ;
        RECT 1.16 2.905 2.805 3.075 ;
        RECT 2.635 2.32 2.805 3.075 ;
        RECT 1.16 2.045 1.33 3.075 ;
        RECT 0.805 2.045 1.33 2.265 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2893 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.47 0.65 0.7 ;
        RECT 0.085 2.435 0.47 3.045 ;
        RECT 0.085 0.47 0.355 3.045 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.735 -0.085 3.065 0.985 ;
        RECT 0.83 -0.085 1.16 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.975 2.66 3.175 3.415 ;
        RECT 0.64 2.435 0.99 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.345 2.66 3.735 2.94 ;
      RECT 3.565 1.035 3.735 2.94 ;
      RECT 2.635 1.175 2.815 1.845 ;
      RECT 2.635 1.175 3.735 1.345 ;
      RECT 3.235 0.795 3.565 1.345 ;
      RECT 1.565 1.815 1.895 2.735 ;
      RECT 1.565 1.815 2.115 1.985 ;
      RECT 1.945 0.67 2.115 1.985 ;
      RECT 0.525 0.87 0.78 1.67 ;
      RECT 0.525 0.87 2.115 1.04 ;
      RECT 1.845 0.67 2.115 1.04 ;
  END
END scs130lp_mux2_0

MACRO scs130lp_mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.49 1.9 2.58 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.46 0.255 2.735 2.615 ;
        RECT 1.54 0.255 2.735 0.535 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.72 3.85 2.13 ;
        RECT 1.19 2.885 3.075 3.055 ;
        RECT 2.905 1.72 3.075 3.055 ;
        RECT 1.19 1.34 1.36 3.055 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.255 0.47 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 2.905 -0.085 3.495 1.035 ;
        RECT 0.65 -0.085 0.98 0.82 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.245 2.3 3.475 3.415 ;
        RECT 0.71 1.815 1.02 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.645 2.3 4.2 2.57 ;
      RECT 4.03 1.38 4.2 2.57 ;
      RECT 3.665 0.705 4.06 1.55 ;
      RECT 2.98 1.22 4.06 1.55 ;
      RECT 2.07 0.99 2.29 2.54 ;
      RECT 0.64 0.99 0.9 1.52 ;
      RECT 0.64 0.99 2.29 1.16 ;
      RECT 1.775 0.705 2.105 1.16 ;
  END
END scs130lp_mux2_1

MACRO scs130lp_mux2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.965 1.55 2.65 2.005 ;
        RECT 1.965 0.935 2.135 2.005 ;
        RECT 1.805 0.935 2.135 1.185 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.36 0.47 2.735 1.38 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.955 0.785 3.275 1.85 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.58 0.255 0.835 1.095 ;
        RECT 0.58 1.85 0.805 3.075 ;
        RECT 0.58 0.255 0.75 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.905 -0.085 3.235 0.615 ;
        RECT 1.045 -0.085 1.375 0.425 ;
        RECT 0.125 -0.085 0.41 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.985 2.515 3.315 3.415 ;
        RECT 0.985 2.855 1.315 3.415 ;
        RECT 0.125 1.815 0.41 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.485 0.275 3.745 2.895 ;
      RECT 1.42 2.175 3.745 2.345 ;
      RECT 3.445 0.275 3.745 2.345 ;
      RECT 1.42 1.395 1.75 2.345 ;
      RECT 2.085 2.515 2.415 2.845 ;
      RECT 1.005 2.515 2.415 2.685 ;
      RECT 1.005 0.595 1.175 2.685 ;
      RECT 0.93 1.275 1.175 1.605 ;
      RECT 1.005 0.595 2.19 0.765 ;
      RECT 1.93 0.255 2.19 0.765 ;
  END
END scs130lp_mux2_2

MACRO scs130lp_mux2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 0.345 1.905 1.525 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.2 2.725 1.525 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.43 1.695 3.255 1.865 ;
        RECT 2.905 1.2 3.255 1.865 ;
        RECT 0.43 1.335 0.69 1.865 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.855 1.755 5.66 1.925 ;
        RECT 5.46 0.39 5.66 1.925 ;
        RECT 3.765 1.065 5.66 1.235 ;
        RECT 5.435 0.39 5.66 1.235 ;
        RECT 4.715 1.755 4.895 3.075 ;
        RECT 4.645 0.255 4.87 1.235 ;
        RECT 3.855 1.755 4.045 3.075 ;
        RECT 3.765 0.255 3.975 1.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 5.04 -0.085 5.265 0.895 ;
        RECT 4.145 -0.085 4.475 0.895 ;
        RECT 2.875 -0.085 3.595 0.69 ;
        RECT 0.87 -0.085 1.33 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.075 2.095 5.405 3.415 ;
        RECT 4.215 2.095 4.545 3.415 ;
        RECT 3.355 2.445 3.685 3.415 ;
        RECT 0.595 2.035 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.975 2.035 2.305 2.335 ;
      RECT 1.975 2.035 3.65 2.215 ;
      RECT 3.425 1.405 3.65 2.215 ;
      RECT 3.425 1.405 5.28 1.585 ;
      RECT 3.425 0.86 3.595 2.215 ;
      RECT 2.085 0.86 3.595 1.03 ;
      RECT 2.085 0.255 2.53 1.03 ;
      RECT 2.925 2.385 3.185 3.075 ;
      RECT 1.545 2.035 1.795 2.735 ;
      RECT 1.545 2.505 3.185 2.675 ;
      RECT 1.545 2.035 1.805 2.675 ;
      RECT 1.095 2.905 2.735 3.075 ;
      RECT 2.405 2.845 2.735 3.075 ;
      RECT 1.095 2.035 1.355 3.075 ;
      RECT 0.09 2.035 0.425 3.075 ;
      RECT 0.09 0.255 0.26 3.075 ;
      RECT 1.085 0.985 1.415 1.525 ;
      RECT 0.09 0.985 1.415 1.155 ;
      RECT 0.09 0.255 0.7 1.155 ;
  END
END scs130lp_mux2_4

MACRO scs130lp_mux2_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_8 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.492 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.765 1.025 7.095 1.395 ;
        RECT 4.975 1.025 7.095 1.195 ;
        RECT 4.815 1.565 5.145 1.895 ;
        RECT 4.975 1.025 5.145 1.895 ;
    END
  END A0
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 0.925 3.525 1.095 ;
        RECT 3.195 0.295 3.525 1.095 ;
        RECT 3.125 1.815 3.375 3.075 ;
        RECT 0.545 1.815 3.375 1.985 ;
        RECT 2.265 1.815 2.595 3.075 ;
        RECT 2.265 0.295 2.595 1.095 ;
        RECT 1.405 1.815 1.735 3.075 ;
        RECT 1.405 0.295 1.735 1.095 ;
        RECT 0.545 0.295 0.875 3.075 ;
    END
  END X
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.192 LAYER li ;
      ANTENNAGATEAREA 0.492 LAYER met1 ;
      ANTENNAMAXAREACAR 0.94349 LAYER li ;
      ANTENNAMAXAREACAR 0.94349 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.130208 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.130208 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.150521 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 6.335 1.55 6.625 1.78 ;
        RECT 4.415 1.595 6.625 1.735 ;
        RECT 4.415 1.55 4.705 1.78 ;
      LAYER li ;
        RECT 6.355 1.565 7.095 1.925 ;
        RECT 6.355 1.55 6.595 1.925 ;
        RECT 4.475 1.025 4.805 1.355 ;
        RECT 4.475 1.025 4.645 1.78 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
      ANTENNAGATEAREA 0.807 LAYER met1 ;
      ANTENNAMAXAREACAR 1.224898 LAYER li ;
      ANTENNAMAXAREACAR 1.224898 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.162602 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.162602 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.091746 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.92 8.065 2.15 ;
        RECT 5.375 1.965 8.065 2.105 ;
        RECT 5.375 1.92 5.665 2.15 ;
      LAYER li ;
        RECT 7.865 1.345 8.37 1.675 ;
        RECT 7.805 1.92 8.035 2.15 ;
        RECT 7.865 1.345 8.035 2.15 ;
        RECT 4.395 2.065 5.685 2.235 ;
        RECT 5.355 1.555 5.685 2.235 ;
        RECT 3.965 1.98 4.565 2.15 ;
        RECT 3.965 1.605 4.305 2.15 ;
    END
  END S
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.64 0.085 ;
        RECT 7.665 -0.085 7.995 0.835 ;
        RECT 5.68 -0.085 6.01 0.515 ;
        RECT 3.705 -0.085 3.955 1.095 ;
        RECT 2.775 -0.085 3.025 0.755 ;
        RECT 1.915 -0.085 2.085 0.755 ;
        RECT 1.055 -0.085 1.225 0.755 ;
        RECT 0.115 -0.085 0.375 1.115 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.64 3.415 ;
        RECT 7.745 2.66 8.075 3.415 ;
        RECT 5.69 2.775 6.02 3.415 ;
        RECT 3.555 2.66 3.885 3.415 ;
        RECT 2.775 2.155 2.945 3.415 ;
        RECT 1.915 2.155 2.085 3.415 ;
        RECT 1.055 2.155 1.225 3.415 ;
        RECT 0.115 1.795 0.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.255 1.845 8.505 3.075 ;
      RECT 7.365 2.32 8.505 2.49 ;
      RECT 7.365 1.005 7.535 2.49 ;
      RECT 6.03 2.095 7.535 2.265 ;
      RECT 5.895 1.555 6.185 2.235 ;
      RECT 7.365 1.005 7.695 1.515 ;
      RECT 7.365 1.005 8.495 1.175 ;
      RECT 8.165 0.255 8.495 1.175 ;
      RECT 6.19 2.905 7.52 3.075 ;
      RECT 7.19 2.66 7.52 3.075 ;
      RECT 6.19 2.775 6.52 3.075 ;
      RECT 7.12 0.295 7.45 0.835 ;
      RECT 6.19 0.295 7.45 0.465 ;
      RECT 6.69 2.435 7.02 2.735 ;
      RECT 4.69 2.405 5.02 2.735 ;
      RECT 5.69 2.435 7.02 2.605 ;
      RECT 4.055 2.405 5.86 2.575 ;
      RECT 3.625 2.32 4.225 2.49 ;
      RECT 3.625 1.265 3.795 2.49 ;
      RECT 1.12 1.265 3.795 1.595 ;
      RECT 1.12 1.265 4.305 1.435 ;
      RECT 4.135 0.685 4.305 1.435 ;
      RECT 4.135 0.685 6.95 0.855 ;
      RECT 6.62 0.635 6.95 0.855 ;
      RECT 4.67 0.595 5 0.855 ;
      RECT 4.19 2.905 5.52 3.075 ;
      RECT 5.19 2.745 5.52 3.075 ;
      RECT 4.19 2.745 4.52 3.075 ;
      RECT 5.17 0.255 5.5 0.515 ;
      RECT 4.17 0.255 4.5 0.515 ;
      RECT 4.17 0.255 5.5 0.425 ;
  END
END scs130lp_mux2_8

MACRO scs130lp_mux2_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.04 1.535 3.235 1.865 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 1.195 2.73 1.365 ;
        RECT 2.4 0.965 2.73 1.365 ;
        RECT 1.5 1.195 1.83 1.78 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.405 1.18 3.735 1.865 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 2.615 0.49 3.075 ;
        RECT 0.115 0.255 0.445 0.715 ;
        RECT 0.115 0.255 0.355 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.065 -0.085 3.395 0.715 ;
        RECT 0.905 -0.085 1.235 0.685 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.59 2.615 2.92 3.415 ;
        RECT 0.95 2.715 1.28 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.845 2.035 4.185 3.075 ;
      RECT 4.015 0.255 4.185 3.075 ;
      RECT 1 2.035 4.185 2.205 ;
      RECT 1 1.835 1.33 2.205 ;
      RECT 3.855 0.255 4.185 0.715 ;
      RECT 1.77 2.375 2.1 3.075 ;
      RECT 0.66 2.375 2.1 2.545 ;
      RECT 0.66 0.885 0.83 2.545 ;
      RECT 0.525 0.885 0.855 1.555 ;
      RECT 1.9 0.255 2.23 1.025 ;
      RECT 0.685 0.855 2.23 1.025 ;
  END
END scs130lp_mux2_lp

MACRO scs130lp_mux2_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_lp2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.985 0.81 2.315 1.145 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.495 0.905 3.235 1.235 ;
        RECT 3.005 0.44 3.235 1.235 ;
        RECT 1.77 1.515 2.665 1.845 ;
        RECT 2.495 0.905 2.665 1.845 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.845 1.475 4.195 1.805 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 0.265 0.45 2.52 ;
        RECT 0.115 0.265 0.445 3.025 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.425 -0.085 3.755 0.725 ;
        RECT 0.91 -0.085 1.24 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.055 2.765 3.385 3.415 ;
        RECT 0.645 2.765 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.585 1.985 3.915 3.025 ;
      RECT 0.91 2.415 3.915 2.585 ;
      RECT 0.91 1.515 1.24 2.585 ;
      RECT 3.585 1.985 4.545 2.155 ;
      RECT 4.375 0.265 4.545 2.155 ;
      RECT 4.215 0.265 4.545 0.725 ;
      RECT 1.42 2.065 2.325 2.235 ;
      RECT 1.42 0.345 1.59 2.235 ;
      RECT 0.63 0.905 1.59 1.235 ;
      RECT 2.495 0.345 2.825 0.725 ;
      RECT 1.42 0.345 2.825 0.515 ;
  END
END scs130lp_mux2_lp2

MACRO scs130lp_mux2_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.445 1.765 1.775 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.295 1.835 2.725 2.165 ;
        RECT 2.295 0.265 2.465 2.165 ;
        RECT 1.515 0.265 2.465 0.435 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 1.58 3.365 2.49 ;
        RECT 2.49 2.345 3.205 2.515 ;
        RECT 1.45 2.895 2.66 3.065 ;
        RECT 2.49 2.345 2.66 3.065 ;
        RECT 1.45 2.015 1.62 3.065 ;
        RECT 1.365 2.015 1.62 2.345 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.231 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.53 0.76 2.86 ;
        RECT 0.155 0.585 0.61 0.915 ;
        RECT 0.155 0.585 0.325 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.645 -0.085 2.975 0.875 ;
        RECT 0.79 -0.085 1.12 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.88 2.695 3.21 3.415 ;
        RECT 0.94 2.675 1.27 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.39 2.67 3.72 2.88 ;
      RECT 3.55 1.155 3.72 2.88 ;
      RECT 2.655 1.155 2.825 1.485 ;
      RECT 2.655 1.155 3.72 1.325 ;
      RECT 3.24 0.795 3.57 1.325 ;
      RECT 1.945 2.525 2.31 2.715 ;
      RECT 1.945 1.095 2.115 2.715 ;
      RECT 0.695 1.095 0.865 2.015 ;
      RECT 0.695 1.095 2.115 1.265 ;
      RECT 1.64 0.795 1.97 1.265 ;
  END
END scs130lp_mux2_m

MACRO scs130lp_mux2i_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2i_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 0.81 2.36 1.985 ;
        RECT 1.46 0.81 2.36 1.38 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 1.55 1.86 1.84 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.385 2.505 3.14 2.675 ;
        RECT 2.87 1.625 3.14 2.675 ;
        RECT 1.47 2.905 2.555 3.075 ;
        RECT 2.385 2.505 2.555 3.075 ;
        RECT 1.47 2.01 1.67 3.075 ;
        RECT 0.535 2.01 1.67 2.245 ;
        RECT 0.535 1.53 0.89 2.245 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4036 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.84 2.165 2.7 2.335 ;
        RECT 2.53 0.285 2.7 2.335 ;
        RECT 1.66 0.285 2.7 0.64 ;
        RECT 1.84 2.165 2.17 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.87 -0.085 3.135 0.615 ;
        RECT 0.705 -0.085 1.035 0.615 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.725 2.845 3.055 3.415 ;
        RECT 0.9 2.435 1.23 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 2.415 0.705 3.055 ;
      RECT 0.085 0.265 0.365 3.055 ;
      RECT 0.085 0.785 1.22 1.36 ;
      RECT 0.085 0.265 0.525 1.36 ;
  END
END scs130lp_mux2i_0

MACRO scs130lp_mux2i_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2i_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.345 0.47 1.76 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.98 1.425 1.31 1.75 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.375 1.21 3.755 1.75 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.693 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.64 1.93 1.285 2.14 ;
        RECT 0.555 0.595 0.885 1.165 ;
        RECT 0.64 0.595 0.81 2.14 ;
        RECT 0.555 0.595 0.81 1.175 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.415 -0.085 3.745 1.04 ;
        RECT 2.085 -0.085 2.305 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.375 1.92 3.705 3.415 ;
        RECT 1.795 2.155 2.125 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.945 1.415 3.205 3.075 ;
      RECT 2.985 0.36 3.205 3.075 ;
      RECT 1.52 1.415 3.205 1.585 ;
      RECT 2.985 0.36 3.245 1.095 ;
      RECT 1.055 1.075 2.775 1.245 ;
      RECT 2.49 0.255 2.775 1.245 ;
      RECT 1.055 0.595 1.385 1.245 ;
      RECT 2.295 1.815 2.595 3.075 ;
      RECT 0.2 2.31 0.53 3.075 ;
      RECT 0.2 2.31 1.625 2.55 ;
      RECT 1.455 1.84 1.625 2.55 ;
      RECT 0.2 1.93 0.47 3.075 ;
      RECT 1.47 1.815 2.595 1.985 ;
      RECT 0.105 0.255 0.385 1.175 ;
      RECT 1.585 0.255 1.915 0.905 ;
      RECT 0.105 0.255 1.915 0.425 ;
  END
END scs130lp_mux2i_1

MACRO scs130lp_mux2i_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2i_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.935 1.425 4.715 1.75 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.885 1.425 5.67 1.75 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.945 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.68 1.405 2.275 1.67 ;
        RECT 0.61 1.855 1.85 2.12 ;
        RECT 1.68 1.405 1.85 2.12 ;
        RECT 0.61 1.345 0.79 2.12 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.785 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.38 1.075 5.59 1.245 ;
        RECT 5.33 0.33 5.59 1.245 ;
        RECT 5.135 1.92 5.43 3.075 ;
        RECT 4.24 1.92 5.43 2.1 ;
        RECT 3.38 0.965 4.65 1.245 ;
        RECT 4.32 0.605 4.65 1.245 ;
        RECT 4.24 1.92 4.57 2.735 ;
        RECT 2.87 1.92 5.43 2.09 ;
        RECT 2.87 1.58 3.71 2.09 ;
        RECT 3.38 0.965 3.71 2.09 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 1.7 0.675 2.85 0.895 ;
        RECT 1.7 -0.085 1.92 0.895 ;
        RECT 0.8 -0.085 1.13 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 2.795 2.94 3.125 3.415 ;
        RECT 1.74 2.94 2.07 3.415 ;
        RECT 0.71 2.29 1.04 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.83 0.255 5.16 0.905 ;
      RECT 2.09 0.255 2.42 0.505 ;
      RECT 2.09 0.255 5.16 0.435 ;
      RECT 3.305 2.905 4.965 3.075 ;
      RECT 4.74 2.27 4.965 3.075 ;
      RECT 1.23 2.29 1.56 2.97 ;
      RECT 3.305 2.6 3.475 3.075 ;
      RECT 1.23 2.6 3.475 2.77 ;
      RECT 1.3 1.065 3.21 1.235 ;
      RECT 3.02 0.605 3.21 1.235 ;
      RECT 1.3 0.255 1.53 1.235 ;
      RECT 3.02 0.605 4.14 0.795 ;
      RECT 3.81 2.26 4.07 2.735 ;
      RECT 2.25 2.26 4.07 2.43 ;
      RECT 2.25 1.84 2.58 2.43 ;
      RECT 0.18 0.255 0.44 3.075 ;
      RECT 0.96 1.415 1.435 1.585 ;
      RECT 0.96 0.985 1.13 1.585 ;
      RECT 0.18 0.985 1.13 1.155 ;
      RECT 0.18 0.255 0.63 1.155 ;
  END
END scs130lp_mux2i_2

MACRO scs130lp_mux2i_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2i_4 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.425 1.715 1.75 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.335 3.775 1.76 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.575 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.855 1.335 9.17 1.665 ;
        RECT 6.875 1.775 9.025 1.945 ;
        RECT 8.855 1.335 9.025 1.945 ;
        RECT 4.435 1.415 7.045 1.835 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.961 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.93 4.265 2.11 ;
        RECT 4.095 0.965 4.265 2.11 ;
        RECT 1.035 0.965 4.265 1.165 ;
        RECT 1.895 0.965 2.255 1.47 ;
        RECT 0.155 1.075 2.255 1.245 ;
        RECT 1.035 0.635 1.365 1.245 ;
        RECT 1.115 1.93 1.285 2.6 ;
        RECT 0.235 1.93 4.265 2.1 ;
        RECT 0.235 1.93 0.425 2.94 ;
        RECT 0.155 0.325 0.345 1.245 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 8.505 -0.085 8.835 0.815 ;
        RECT 7.645 -0.085 7.975 0.805 ;
        RECT 6.855 -0.085 7.115 0.905 ;
        RECT 5.995 -0.085 6.185 0.565 ;
        RECT 5.135 -0.085 5.325 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 8.745 2.125 9.025 3.415 ;
        RECT 7.735 2.455 8.065 3.415 ;
        RECT 6.795 2.845 7.125 3.415 ;
        RECT 5.915 2.845 6.245 3.415 ;
        RECT 4.94 2.97 5.27 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.195 1.845 9.51 3.075 ;
      RECT 9.34 0.985 9.51 3.075 ;
      RECT 7.225 1.415 8.675 1.605 ;
      RECT 8.505 0.985 8.675 1.605 ;
      RECT 8.505 0.985 9.51 1.165 ;
      RECT 9.005 0.255 9.205 1.165 ;
      RECT 2.385 2.63 3.455 3.075 ;
      RECT 8.235 2.115 8.575 3.065 ;
      RECT 7.295 2.115 7.565 3.065 ;
      RECT 2.385 2.63 4.965 2.8 ;
      RECT 6.88 2.115 7.565 2.675 ;
      RECT 4.795 2.505 7.565 2.675 ;
      RECT 6.88 2.115 8.575 2.285 ;
      RECT 4.445 1.075 8.335 1.245 ;
      RECT 8.145 0.255 8.335 1.245 ;
      RECT 7.285 0.255 7.475 1.245 ;
      RECT 4.445 0.625 4.615 1.245 ;
      RECT 0.525 0.255 0.855 0.905 ;
      RECT 1.535 0.625 4.615 0.795 ;
      RECT 1.535 0.255 1.795 0.795 ;
      RECT 0.525 0.255 1.795 0.455 ;
      RECT 4.795 0.735 6.685 0.905 ;
      RECT 6.355 0.255 6.685 0.905 ;
      RECT 5.495 0.345 5.825 0.905 ;
      RECT 4.795 0.255 4.965 0.905 ;
      RECT 2.405 0.255 4.965 0.455 ;
      RECT 0.665 2.78 1.735 2.95 ;
      RECT 1.525 2.28 1.735 2.95 ;
      RECT 0.665 2.28 0.875 2.95 ;
      RECT 1.525 2.28 4.615 2.46 ;
      RECT 4.445 2.005 6.615 2.335 ;
  END
END scs130lp_mux2i_4

MACRO scs130lp_mux2i_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2i_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.725 0.865 2.15 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 2.115 1.585 2.445 ;
        RECT 1.035 1.155 1.205 2.445 ;
        RECT 0.605 1.155 1.205 1.485 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.72 0.775 2.725 1.105 ;
        RECT 1.72 0.255 1.89 1.105 ;
        RECT 0.615 0.255 1.89 0.425 ;
        RECT 0.105 0.815 0.785 0.985 ;
        RECT 0.615 0.255 0.785 0.985 ;
        RECT 0.105 0.815 0.435 1.485 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4014 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.755 1.775 2.275 2.615 ;
        RECT 0.99 2.615 1.925 2.785 ;
        RECT 1.38 1.775 2.275 1.945 ;
        RECT 1.38 0.595 1.55 1.945 ;
        RECT 1.05 0.595 1.55 0.925 ;
        RECT 0.99 2.615 1.32 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.06 -0.085 2.39 0.605 ;
        RECT 0.115 -0.085 0.445 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.095 2.785 2.425 3.415 ;
        RECT 0.17 2.615 0.5 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.885 1.275 3.24 3.075 ;
      RECT 2.91 0.255 3.24 3.075 ;
      RECT 1.825 1.275 3.24 1.605 ;
  END
END scs130lp_mux2i_lp

MACRO scs130lp_mux2i_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2i_lp2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.065 2.24 1.395 ;
        RECT 0.98 1.465 1.73 1.795 ;
        RECT 1.56 1.065 1.73 1.795 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.91 1.605 2.275 2.15 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.715 3.2 1.095 ;
        RECT 1.21 0.715 3.2 0.885 ;
        RECT 0.44 1.075 1.38 1.245 ;
        RECT 1.21 0.715 1.38 1.245 ;
        RECT 0.44 1.075 0.77 1.745 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6918 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.86 0.265 1.98 0.535 ;
        RECT 0.605 2.895 1.825 3.065 ;
        RECT 1.495 2.33 1.825 3.065 ;
        RECT 0.605 2.095 1.315 3.065 ;
        RECT 0.09 0.725 1.03 0.895 ;
        RECT 0.86 0.265 1.03 0.895 ;
        RECT 0.09 1.925 0.775 2.095 ;
        RECT 0.09 0.725 0.26 2.095 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.58 -0.085 2.91 0.535 ;
        RECT 0.35 -0.085 0.68 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.705 2.075 3.035 3.415 ;
        RECT 0.175 2.275 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.275 1.335 3.71 3.065 ;
      RECT 3.38 0.265 3.71 3.065 ;
      RECT 2.48 1.335 3.71 1.665 ;
  END
END scs130lp_mux2i_lp2

MACRO scs130lp_mux2i_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux2i_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 1.58 2.36 1.795 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.355 0.265 2.15 0.435 ;
        RECT 1.355 1.21 1.765 2.12 ;
        RECT 1.355 0.265 1.525 2.12 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.295 2.325 3.205 2.495 ;
        RECT 2.89 1.155 3.205 2.495 ;
        RECT 1.335 2.895 2.465 3.065 ;
        RECT 2.295 2.325 2.465 3.065 ;
        RECT 1.335 2.3 1.505 3.065 ;
        RECT 0.52 2.3 1.505 2.47 ;
        RECT 0.52 1.995 0.69 2.47 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 1.975 2.71 2.145 ;
        RECT 2.54 1.055 2.71 2.145 ;
        RECT 2.075 1.055 2.71 1.225 ;
        RECT 2.075 0.7 2.245 1.225 ;
        RECT 1.71 2.525 2.115 2.715 ;
        RECT 1.945 1.975 2.115 2.715 ;
        RECT 1.705 0.7 2.245 1.03 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.6 -0.085 2.93 0.875 ;
        RECT 0.745 -0.085 1.075 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.79 2.675 3.12 3.415 ;
        RECT 0.825 2.655 1.155 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.17 2.65 0.645 2.86 ;
      RECT 0.17 0.795 0.34 2.86 ;
      RECT 0.17 1.425 1.17 1.755 ;
      RECT 0.17 0.795 0.565 1.005 ;
  END
END scs130lp_mux2i_m

MACRO scs130lp_mux4_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux4_0 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.215 1.14 4.725 1.39 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 1.145 3.685 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.55 1.93 1.11 2.19 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.34 1.93 2.845 2.13 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.29 1.94 1.68 2.19 ;
        RECT 1.29 1.58 1.46 2.19 ;
        RECT 0.47 1.375 1.29 1.76 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.66 0.78 7.115 1.825 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.285 0.28 7.585 2.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.86 -0.085 7.115 0.61 ;
        RECT 4.335 -0.085 4.665 0.97 ;
        RECT 2.655 -0.085 2.985 0.97 ;
        RECT 0.895 -0.085 1.225 0.865 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.915 1.995 7.095 3.415 ;
        RECT 6.88 1.995 7.095 2.675 ;
        RECT 6.8 1.995 7.095 2.615 ;
        RECT 4.3 2.67 4.63 3.415 ;
        RECT 2.67 2.64 2.92 3.415 ;
        RECT 0.615 2.7 0.945 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 5.855 0.81 6.145 1.04 ;
      RECT 2.015 0.81 2.305 1.04 ;
      RECT 2.015 0.855 6.145 0.995 ;
    LAYER li ;
      RECT 5.42 2.905 6.745 3.075 ;
      RECT 6.415 2.78 6.745 3.075 ;
      RECT 5.42 0.67 5.61 3.075 ;
      RECT 5.42 0.67 5.64 1.005 ;
      RECT 6.3 2.06 6.63 2.39 ;
      RECT 6.3 1.525 6.49 2.39 ;
      RECT 6.31 0.255 6.49 2.39 ;
      RECT 6.12 1.525 6.49 1.855 ;
      RECT 6.31 0.255 6.69 0.61 ;
      RECT 5.145 0.255 6.69 0.5 ;
      RECT 5.78 2.46 6.11 2.735 ;
      RECT 5.78 1.175 5.95 2.735 ;
      RECT 5.81 0.67 6.14 1.345 ;
      RECT 3.455 2.64 3.875 2.92 ;
      RECT 3.705 2.33 3.875 2.92 ;
      RECT 4.92 2.33 5.25 2.84 ;
      RECT 5.08 0.67 5.25 2.84 ;
      RECT 3.705 2.33 5.25 2.5 ;
      RECT 3.865 1.56 5.25 1.73 ;
      RECT 4.95 0.67 5.25 1.73 ;
      RECT 3.865 0.64 4.035 1.73 ;
      RECT 3.545 0.64 4.035 0.97 ;
      RECT 1.135 2.905 2.5 3.075 ;
      RECT 2.33 2.3 2.5 3.075 ;
      RECT 0.115 2.36 0.445 2.905 ;
      RECT 1.135 2.36 1.305 3.075 ;
      RECT 0.115 2.36 1.305 2.53 ;
      RECT 2.33 2.3 3.535 2.47 ;
      RECT 3.275 1.93 3.535 2.47 ;
      RECT 0.115 1.025 0.3 2.905 ;
      RECT 3.275 1.93 4.9 2.16 ;
      RECT 1.63 1.195 1.82 1.685 ;
      RECT 1.485 1.195 1.82 1.365 ;
      RECT 0.115 1.035 1.655 1.205 ;
      RECT 0.115 1.025 0.725 1.205 ;
      RECT 0.465 0.64 0.725 1.205 ;
      RECT 1.56 2.475 2.16 2.735 ;
      RECT 1.99 0.64 2.16 2.735 ;
      RECT 1.99 0.64 2.325 1.015 ;
      RECT 1.825 0.64 2.325 0.97 ;
  END
END scs130lp_mux4_0

MACRO scs130lp_mux4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux4_1 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.83 1.175 1.45 2.175 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.155 0.55 2.175 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.4 1.21 5.88 1.765 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.945 1.08 5.23 1.765 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.99 1.125 3.65 1.795 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.795 1.355 7.125 1.865 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.725 0.375 9.995 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.225 -0.085 9.555 1.175 ;
        RECT 6.49 -0.085 6.82 0.845 ;
        RECT 5.39 -0.085 5.72 0.475 ;
        RECT 2.99 -0.085 3.32 0.955 ;
        RECT 0.555 -0.085 0.885 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.225 1.845 9.555 3.415 ;
        RECT 6.41 2.375 6.75 3.415 ;
        RECT 5.285 2.615 5.535 3.415 ;
        RECT 3.345 2.515 3.645 3.415 ;
        RECT 0.525 2.685 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 7.775 1.92 8.065 2.15 ;
      RECT 2.015 1.92 2.305 2.15 ;
      RECT 2.015 1.965 8.065 2.105 ;
    LAYER li ;
      RECT 8.22 0.79 8.44 2.21 ;
      RECT 8.22 1.345 9.555 1.675 ;
      RECT 8.22 0.79 8.445 1.675 ;
      RECT 7.78 1.88 8.05 2.21 ;
      RECT 7.88 0.39 8.05 2.21 ;
      RECT 8.615 0.39 8.91 1.12 ;
      RECT 7.88 0.39 8.91 0.62 ;
      RECT 4.385 2.525 4.775 2.735 ;
      RECT 4.605 1.015 4.775 2.735 ;
      RECT 7.43 2.38 8.85 2.61 ;
      RECT 8.61 1.88 8.85 2.61 ;
      RECT 7.43 0.79 7.6 2.61 ;
      RECT 6.445 2.035 7.6 2.205 ;
      RECT 4.605 1.935 6.615 2.105 ;
      RECT 3.975 1.015 4.775 1.185 ;
      RECT 7.43 0.79 7.71 1.12 ;
      RECT 3.975 0.625 4.2 1.185 ;
      RECT 6.92 2.78 7.65 3.075 ;
      RECT 6.92 2.375 7.25 3.075 ;
      RECT 6.225 1.015 6.555 1.765 ;
      RECT 6.225 1.015 7.25 1.185 ;
      RECT 7 0.64 7.25 1.185 ;
      RECT 4.37 0.645 6.16 0.845 ;
      RECT 5.89 0.275 6.16 0.845 ;
      RECT 4.37 0.615 4.7 0.845 ;
      RECT 3.955 2.905 5.115 3.075 ;
      RECT 4.945 2.275 5.115 3.075 ;
      RECT 3.955 2.545 4.205 3.075 ;
      RECT 5.705 2.275 6.005 2.88 ;
      RECT 4.945 2.275 6.005 2.445 ;
      RECT 3.51 0.255 3.805 0.955 ;
      RECT 4.89 0.255 5.22 0.475 ;
      RECT 3.51 0.255 5.22 0.445 ;
      RECT 2.885 1.975 3.175 2.845 ;
      RECT 2.65 1.975 4.435 2.145 ;
      RECT 4.175 1.365 4.435 2.145 ;
      RECT 2.65 0.64 2.82 2.145 ;
      RECT 2.255 1.1 2.82 1.77 ;
      RECT 2.56 0.64 2.82 1.77 ;
      RECT 1.025 2.865 2.665 3.035 ;
      RECT 2.405 2.34 2.665 3.035 ;
      RECT 1.025 2.685 1.285 3.035 ;
      RECT 1.905 1.94 2.235 2.67 ;
      RECT 1.905 1.94 2.305 2.17 ;
      RECT 1.905 0.835 2.075 2.67 ;
      RECT 1.395 0.835 2.075 1.005 ;
      RECT 1.395 0.615 1.725 1.005 ;
      RECT 0.125 0.815 1.225 0.985 ;
      RECT 1.055 0.265 1.225 0.985 ;
      RECT 0.125 0.45 0.385 0.985 ;
      RECT 1.895 0.265 2.225 0.665 ;
      RECT 1.055 0.265 2.225 0.435 ;
      RECT 0.095 2.345 0.355 2.97 ;
      RECT 1.475 2.345 1.735 2.675 ;
      RECT 0.095 2.345 1.735 2.515 ;
  END
END scs130lp_mux4_1

MACRO scs130lp_mux4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux4_2 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.685 1.57 7.62 1.855 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.785 1.345 6.165 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.685 1.57 5.615 1.905 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.425 1.145 4.165 2.265 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.477 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.79 1.325 8.12 1.905 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.285 2.325 2.12 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 0.255 3.255 2.265 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.64 0.085 ;
        RECT 7.35 -0.085 7.68 0.815 ;
        RECT 5.485 -0.085 5.815 0.825 ;
        RECT 3.425 -0.085 4.015 0.975 ;
        RECT 2.485 -0.085 2.815 0.355 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.64 3.415 ;
        RECT 7.485 2.085 7.815 3.415 ;
        RECT 5.21 2.29 5.99 3.415 ;
        RECT 5.21 2.075 5.54 3.415 ;
        RECT 3.385 2.785 3.715 3.415 ;
        RECT 2.525 2.785 2.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 6.335 2.29 6.625 2.52 ;
      RECT 1.055 2.29 1.345 2.52 ;
      RECT 1.055 2.335 6.625 2.475 ;
    LAYER li ;
      RECT 7.985 2.075 8.47 2.745 ;
      RECT 8.3 0.985 8.47 2.745 ;
      RECT 6.685 0.985 7.13 1.4 ;
      RECT 6.96 0.265 7.13 1.4 ;
      RECT 4.695 0.995 5.025 1.4 ;
      RECT 4.695 0.995 6.155 1.165 ;
      RECT 5.985 0.265 6.155 1.165 ;
      RECT 6.685 0.985 8.47 1.155 ;
      RECT 7.85 0.64 8.11 1.155 ;
      RECT 5.985 0.265 7.13 0.435 ;
      RECT 6.335 2.075 6.83 2.745 ;
      RECT 6.335 0.605 6.515 2.745 ;
      RECT 6.335 0.605 6.78 0.815 ;
      RECT 0.095 2.815 1.635 2.985 ;
      RECT 1.465 2.435 1.635 2.985 ;
      RECT 0.095 0.67 0.385 2.985 ;
      RECT 4.42 2.075 4.75 2.745 ;
      RECT 1.465 2.435 4.75 2.605 ;
      RECT 4.345 0.565 4.515 2.605 ;
      RECT 4.345 0.565 4.79 0.825 ;
      RECT 0.555 0.325 0.775 2.635 ;
      RECT 2.605 0.525 2.855 1.515 ;
      RECT 1.465 0.525 2.855 0.695 ;
      RECT 1.465 0.325 1.635 0.695 ;
      RECT 0.555 0.325 1.635 0.495 ;
      RECT 1.565 1.065 1.895 2.265 ;
      RECT 1.295 1.065 1.895 1.825 ;
      RECT 1.725 0.865 2.155 1.115 ;
      RECT 0.955 1.995 1.295 2.575 ;
      RECT 0.955 0.665 1.125 2.575 ;
      RECT 0.955 0.665 1.285 0.895 ;
  END
END scs130lp_mux4_2

MACRO scs130lp_mux4_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux4_4 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.225 1.58 6.565 1.91 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.475 1.185 4.68 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.835 1.485 8.265 2.86 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.765 1.58 7.045 1.91 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.477 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.795 0.47 8.985 1.795 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.185 2.245 2.12 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.865 1.21 4.165 1.815 ;
        RECT 3.865 0.36 4.035 1.815 ;
        RECT 2.815 1.645 3.865 1.985 ;
        RECT 2.965 0.86 4.035 1.03 ;
        RECT 3.825 0.36 4.035 1.03 ;
        RECT 2.965 0.36 3.175 1.03 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 8.07 -0.085 8.4 0.845 ;
        RECT 5.965 -0.085 6.295 0.7 ;
        RECT 4.255 -0.085 4.465 0.885 ;
        RECT 3.395 -0.085 3.605 0.545 ;
        RECT 2.555 -0.085 2.745 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 8.49 2.425 8.7 3.415 ;
        RECT 6.27 2.485 6.6 3.415 ;
        RECT 4.395 2.345 4.725 3.415 ;
        RECT 3.185 2.725 3.515 3.415 ;
        RECT 2.325 2.725 2.655 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 7.295 0.44 7.585 0.67 ;
      RECT 0.095 0.44 0.385 0.67 ;
      RECT 0.095 0.485 7.585 0.625 ;
    LAYER li ;
      RECT 8.92 1.975 9.13 2.745 ;
      RECT 8.445 1.975 9.495 2.145 ;
      RECT 9.165 0.765 9.495 2.145 ;
      RECT 8.445 1.125 8.615 2.145 ;
      RECT 5.605 1.485 6.045 1.815 ;
      RECT 5.875 1.23 6.045 1.815 ;
      RECT 7.485 1.125 7.655 1.795 ;
      RECT 5.875 1.23 7.655 1.4 ;
      RECT 7.485 1.125 8.615 1.295 ;
      RECT 7.41 2.09 7.62 2.76 ;
      RECT 5.255 2.09 7.62 2.26 ;
      RECT 5.255 1.135 5.425 2.26 ;
      RECT 5.255 1.135 5.695 1.305 ;
      RECT 5.525 0.88 5.695 1.305 ;
      RECT 5.525 0.88 6.645 1.05 ;
      RECT 7.23 0.47 7.525 0.905 ;
      RECT 6.475 0.735 7.525 0.905 ;
      RECT 4.905 2.44 5.6 2.77 ;
      RECT 1.035 0.64 1.245 2.67 ;
      RECT 1.035 2.37 4.215 2.54 ;
      RECT 4.045 1.995 4.215 2.54 ;
      RECT 4.905 0.625 5.075 2.77 ;
      RECT 4.045 1.995 5.075 2.165 ;
      RECT 4.905 0.625 5.345 0.955 ;
      RECT 0.605 0.29 0.795 2.66 ;
      RECT 2.615 1.265 3.64 1.435 ;
      RECT 2.615 0.835 2.785 1.435 ;
      RECT 2.205 0.835 2.785 1.005 ;
      RECT 2.205 0.29 2.375 1.005 ;
      RECT 0.605 0.29 2.375 0.46 ;
      RECT 1.565 1.15 1.895 2.19 ;
      RECT 1.725 0.64 1.895 2.19 ;
      RECT 1.425 1.15 1.895 1.82 ;
      RECT 1.725 0.64 2.025 0.97 ;
      RECT 0.155 0.47 0.365 2.66 ;
  END
END scs130lp_mux4_4

MACRO scs130lp_mux4_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux4_lp 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.285 1.21 9.475 1.46 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.74 1.08 7.075 1.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.77 0.765 6.085 1.095 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 1.55 4.35 2.15 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.002 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.18 1.64 9.62 2.15 ;
        RECT 7.44 2.545 8.35 2.715 ;
        RECT 8.18 1.64 8.35 2.715 ;
        RECT 7.44 1.08 7.61 2.715 ;
        RECT 6.325 1.59 7.61 1.76 ;
        RECT 7.28 1.08 7.61 1.76 ;
        RECT 6.325 1.275 6.495 1.76 ;
        RECT 5.395 1.275 6.495 1.445 ;
        RECT 5.815 1.275 6.145 1.76 ;
        RECT 4.885 1.045 5.565 1.375 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.335 1.55 2.755 1.89 ;
        RECT 1.635 2.545 2.505 2.715 ;
        RECT 2.335 1.55 2.505 2.715 ;
        RECT 1.635 1.47 1.805 2.715 ;
        RECT 1.03 1.47 1.805 1.8 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 0.265 0.445 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.845 -0.085 9.175 0.675 ;
        RECT 6.615 -0.085 6.865 0.55 ;
        RECT 3.755 -0.085 4.005 0.945 ;
        RECT 0.905 -0.085 1.235 0.465 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.985 2.68 9.315 3.415 ;
        RECT 6.58 2.29 6.91 3.415 ;
        RECT 3.855 2.865 4.185 3.415 ;
        RECT 0.645 2.33 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.515 2.33 9.97 3.065 ;
      RECT 9.8 0.265 9.97 3.065 ;
      RECT 7.09 2.895 8.805 3.065 ;
      RECT 8.635 2.33 8.805 3.065 ;
      RECT 7.09 1.94 7.26 3.065 ;
      RECT 8.635 2.33 9.97 2.5 ;
      RECT 5.465 1.94 7.26 2.11 ;
      RECT 5.465 1.745 5.635 2.11 ;
      RECT 4.885 1.745 5.635 1.915 ;
      RECT 4.885 1.585 5.215 1.915 ;
      RECT 8.14 0.86 9.97 1.03 ;
      RECT 9.635 0.265 9.97 1.03 ;
      RECT 8.14 0.765 8.47 1.03 ;
      RECT 2.685 2.165 2.935 2.715 ;
      RECT 7.79 0.265 7.96 2.365 ;
      RECT 2.685 2.165 3.765 2.335 ;
      RECT 3.595 1.125 3.765 2.335 ;
      RECT 3.395 1.125 4.355 1.295 ;
      RECT 4.185 0.265 4.355 1.295 ;
      RECT 3.395 0.265 3.565 1.295 ;
      RECT 6.265 0.73 7.96 0.9 ;
      RECT 7.545 0.265 7.96 0.9 ;
      RECT 6.265 0.265 6.435 0.9 ;
      RECT 2.325 0.265 2.655 0.725 ;
      RECT 4.185 0.265 6.435 0.435 ;
      RECT 2.325 0.265 3.565 0.435 ;
      RECT 4.955 2.095 5.285 3.065 ;
      RECT 1.205 2.895 3.285 3.065 ;
      RECT 3.115 2.515 3.285 3.065 ;
      RECT 1.205 1.98 1.455 3.065 ;
      RECT 3.115 2.515 5.285 2.685 ;
      RECT 4.535 0.615 4.705 2.685 ;
      RECT 0.625 1.98 1.455 2.15 ;
      RECT 0.625 0.645 0.795 2.15 ;
      RECT 4.535 0.615 5.355 0.865 ;
      RECT 0.625 0.645 1.795 0.815 ;
      RECT 1.465 0.265 1.795 0.815 ;
      RECT 3.045 1.655 3.415 1.985 ;
      RECT 3.045 0.615 3.215 1.985 ;
      RECT 2.335 0.99 3.215 1.32 ;
      RECT 2.885 0.615 3.215 1.32 ;
      RECT 1.985 0.995 2.155 2.365 ;
      RECT 0.975 0.995 2.155 1.26 ;
      RECT 1.975 0.265 2.145 1.26 ;
  END
END scs130lp_mux4_lp

MACRO scs130lp_mux4_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_mux4_m 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.315 1.16 4.645 1.49 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.47 3.235 1.98 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.485 1.285 2.86 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.365 1.47 2.725 1.98 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.265 0.675 0.435 ;
        RECT 0.155 0.265 0.325 0.64 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.795 0.84 7.125 1.355 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.795 0.345 8.005 2.945 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.385 -0.085 7.575 0.545 ;
        RECT 4.265 -0.085 4.475 0.94 ;
        RECT 2.705 -0.085 2.895 0.92 ;
        RECT 0.88 -0.085 1.21 0.88 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.365 2.745 7.575 3.415 ;
        RECT 4.575 2.425 4.745 3.415 ;
        RECT 2.495 2.525 2.825 3.415 ;
        RECT 0.745 2.425 0.935 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.975 0.965 6.165 2.625 ;
      RECT 7.445 1.19 7.615 1.86 ;
      RECT 5.975 1.535 7.615 1.705 ;
      RECT 6.935 0.265 7.145 0.595 ;
      RECT 5.59 0.265 7.145 0.435 ;
      RECT 6.935 1.885 7.145 2.945 ;
      RECT 6.345 1.885 7.145 2.055 ;
      RECT 4.925 2.805 6.595 2.975 ;
      RECT 6.385 2.425 6.595 2.975 ;
      RECT 3.005 2.745 4.395 2.915 ;
      RECT 4.225 2.075 4.395 2.915 ;
      RECT 5.625 0.615 5.795 2.975 ;
      RECT 4.925 2.075 5.095 2.975 ;
      RECT 3.005 2.175 3.175 2.915 ;
      RECT 1.76 2.175 2.005 2.625 ;
      RECT 1.76 2.175 3.175 2.345 ;
      RECT 4.225 2.075 5.095 2.245 ;
      RECT 2.005 0.625 2.175 2.345 ;
      RECT 6.385 0.615 6.595 1.165 ;
      RECT 1.87 0.625 2.175 0.955 ;
      RECT 5.625 0.615 6.595 0.785 ;
      RECT 5.275 0.965 5.445 2.625 ;
      RECT 3.57 2.355 4.045 2.565 ;
      RECT 3.875 0.71 4.045 2.565 ;
      RECT 3.875 1.725 5.445 1.895 ;
      RECT 5.255 0.965 5.445 1.895 ;
      RECT 3.415 0.71 4.045 0.92 ;
      RECT 0.315 0.82 0.525 2.625 ;
      RECT 3.525 1.1 3.695 1.88 ;
      RECT 1.52 1.135 1.825 1.83 ;
      RECT 0.315 1.135 1.825 1.305 ;
      RECT 2.355 1.1 3.695 1.27 ;
      RECT 1.52 0.275 1.69 1.83 ;
      RECT 0.315 0.82 0.7 1.305 ;
      RECT 2.355 0.275 2.525 1.27 ;
      RECT 1.52 0.275 2.525 0.445 ;
  END
END scs130lp_mux4_m

MACRO scs130lp_nand2_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_0 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.84 1.355 2.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.435 2.12 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2905 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 0.28 1.315 0.61 ;
        RECT 0.605 0.28 0.815 2.97 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.165 -0.085 0.435 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.985 2.29 1.315 3.415 ;
        RECT 0.125 2.29 0.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand2_0

MACRO scs130lp_nand2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.21 1.355 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.435 1.75 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5754 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 0.36 1.255 1.04 ;
        RECT 0.605 0.36 0.815 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.105 -0.085 0.435 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.985 1.92 1.295 3.415 ;
        RECT 0.105 1.92 0.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand2_1

MACRO scs130lp_nand2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.1 1.415 1.83 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.415 0.93 1.75 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9408 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.92 2.31 2.09 ;
        RECT 2 1.075 2.31 2.09 ;
        RECT 1.385 1.075 2.31 1.245 ;
        RECT 1.385 0.605 1.715 1.245 ;
        RECT 1.455 1.92 1.645 3.075 ;
        RECT 0.595 1.92 0.785 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.525 -0.085 0.855 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.815 2.26 2.145 3.415 ;
        RECT 0.955 2.27 1.285 3.415 ;
        RECT 0.095 1.925 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.095 1.075 1.205 1.245 ;
      RECT 1.035 0.265 1.205 1.245 ;
      RECT 0.095 0.305 0.355 1.245 ;
      RECT 1.895 0.265 2.225 0.895 ;
      RECT 1.035 0.265 2.225 0.435 ;
  END
END scs130lp_nand2_2

MACRO scs130lp_nand2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_4 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.925 1.415 3.77 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.425 2.245 1.76 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8816 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.075 3.775 1.245 ;
        RECT 3.435 0.605 3.775 1.245 ;
        RECT 3.42 1.93 3.77 3.055 ;
        RECT 0.635 1.93 3.77 2.14 ;
        RECT 2.425 0.615 2.755 2.14 ;
        RECT 2.495 0.615 2.75 3.055 ;
        RECT 1.635 1.93 1.825 3.055 ;
        RECT 0.635 1.93 0.965 3.055 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 1.565 -0.085 1.895 0.915 ;
        RECT 0.705 -0.085 1.035 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.94 1.815 4.205 3.415 ;
        RECT 2.92 2.31 3.25 3.415 ;
        RECT 1.995 2.31 2.325 3.415 ;
        RECT 1.135 2.31 1.465 3.415 ;
        RECT 0.125 1.805 0.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.285 1.085 2.255 1.255 ;
      RECT 2.065 0.265 2.255 1.255 ;
      RECT 3.945 0.265 4.205 1.185 ;
      RECT 1.205 0.305 1.395 1.255 ;
      RECT 0.285 0.305 0.535 1.255 ;
      RECT 2.935 0.265 3.265 0.905 ;
      RECT 2.065 0.265 4.205 0.435 ;
  END
END scs130lp_nand2_4

MACRO scs130lp_nand2_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_8 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.43 1.425 5.78 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.815 1.415 3.505 1.605 ;
        RECT 1.815 1.415 2.825 1.76 ;
        RECT 0.455 1.415 3.505 1.595 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.9732 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.785 0.605 7.115 1.5 ;
        RECT 6.855 0.605 7.055 3.075 ;
        RECT 5.95 1.155 7.055 1.925 ;
        RECT 3.965 1.085 6.22 1.255 ;
        RECT 5.965 0.605 6.22 1.925 ;
        RECT 5.95 1.075 6.185 3.075 ;
        RECT 4.035 1.93 6.185 2.1 ;
        RECT 4.965 1.075 6.22 1.255 ;
        RECT 4.965 0.595 5.295 1.255 ;
        RECT 4.93 1.93 5.26 3.075 ;
        RECT 3.965 0.595 4.295 1.255 ;
        RECT 4.035 0.595 4.26 3.075 ;
        RECT 3.965 0.595 4.26 1.945 ;
        RECT 3.125 1.775 4.26 1.945 ;
        RECT 3.175 1.775 3.365 3.075 ;
        RECT 1.455 1.93 3.365 2.1 ;
        RECT 2.315 1.93 2.505 3.075 ;
        RECT 1.455 1.93 1.645 3.075 ;
        RECT 0.595 1.765 1.635 1.935 ;
        RECT 0.595 1.765 0.785 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 3.105 -0.085 3.435 0.905 ;
        RECT 2.245 -0.085 2.575 0.905 ;
        RECT 1.385 -0.085 1.715 0.905 ;
        RECT 0.525 -0.085 0.855 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.275 1.815 7.485 3.415 ;
        RECT 6.355 2.095 6.685 3.415 ;
        RECT 5.43 2.27 5.76 3.415 ;
        RECT 4.43 2.27 4.76 3.415 ;
        RECT 3.535 2.115 3.865 3.415 ;
        RECT 2.675 2.27 3.005 3.415 ;
        RECT 1.815 2.27 2.145 3.415 ;
        RECT 0.955 2.105 1.285 3.415 ;
        RECT 0.095 1.82 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.095 1.075 3.795 1.245 ;
      RECT 3.605 0.255 3.795 1.245 ;
      RECT 7.285 0.255 7.545 1.19 ;
      RECT 2.745 0.305 2.935 1.245 ;
      RECT 1.885 0.305 2.075 1.245 ;
      RECT 1.025 0.305 1.205 1.245 ;
      RECT 0.095 0.305 0.355 1.245 ;
      RECT 6.39 0.255 6.615 0.985 ;
      RECT 4.465 0.255 4.795 0.915 ;
      RECT 5.465 0.255 5.795 0.905 ;
      RECT 5.465 0.255 7.545 0.435 ;
      RECT 3.605 0.255 7.545 0.425 ;
  END
END scs130lp_nand2_8

MACRO scs130lp_nand2_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_lp 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.93 1.18 1.315 1.575 ;
        RECT 0.93 0.905 1.22 1.575 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.955 0.4 2.89 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2373 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.58 1.815 1.315 2.275 ;
        RECT 0.58 0.555 1.3 0.725 ;
        RECT 0.97 0.265 1.3 0.725 ;
        RECT 0.58 0.555 0.75 2.275 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.15 -0.085 0.4 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.58 2.505 0.91 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand2_lp

MACRO scs130lp_nand2_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_lp2 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 0.85 1.325 1.52 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.55 1.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3997 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.73 1.7 1.795 1.87 ;
        RECT 1.625 0.44 1.795 1.87 ;
        RECT 1.085 0.44 1.795 0.67 ;
        RECT 1.085 0.265 1.45 0.67 ;
        RECT 0.73 1.7 1.06 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.3 -0.085 0.63 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.26 2.05 1.59 3.415 ;
        RECT 0.2 2.025 0.53 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand2_lp2

MACRO scs130lp_nand2_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2_m 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.84 1.285 2.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.435 2.12 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.615 0.33 1.255 0.66 ;
        RECT 0.615 0.33 0.805 2.97 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.225 -0.085 0.435 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 1.045 2.3 1.255 3.415 ;
        RECT 0.185 2.3 0.395 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand2_m

MACRO scs130lp_nand2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2b_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.015 0.455 1.525 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.015 1.285 1.435 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6384 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.945 2.315 2.115 ;
        RECT 2.07 0.255 2.315 2.115 ;
        RECT 1.795 0.255 2.315 1.095 ;
        RECT 1.115 1.945 1.375 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.81 -0.085 1.14 0.505 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.545 2.285 1.875 3.415 ;
        RECT 0.685 2.035 0.945 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.16 1.695 0.49 2.21 ;
      RECT 0.16 1.695 0.78 1.865 ;
      RECT 0.61 1.605 1.635 1.775 ;
      RECT 1.455 1.275 1.9 1.605 ;
      RECT 1.455 0.675 1.625 1.775 ;
      RECT 0.38 0.675 1.625 0.845 ;
      RECT 0.38 0.28 0.64 0.845 ;
  END
END scs130lp_nand2b_1

MACRO scs130lp_nand2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2b_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.185 0.84 1.515 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.365 1.075 2.695 1.515 ;
        RECT 1.01 1.075 2.695 1.245 ;
        RECT 1.01 1.075 1.3 1.515 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9702 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.875 0.725 3.275 2.12 ;
        RECT 1.97 1.83 3.275 2.12 ;
        RECT 1.63 0.725 3.275 0.905 ;
        RECT 2.13 1.83 2.32 3.075 ;
        RECT 1.23 2.035 2.32 2.205 ;
        RECT 1.63 0.655 1.96 0.905 ;
        RECT 1.23 2.035 1.46 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.56 -0.085 2.82 0.555 ;
        RECT 0.525 -0.085 0.95 0.905 ;
        RECT 0.525 -0.085 0.855 0.995 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.49 2.29 2.82 3.415 ;
        RECT 1.63 2.375 1.96 3.415 ;
        RECT 0.675 2.035 1.06 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.12 0.255 1.45 0.905 ;
      RECT 1.12 0.255 2.39 0.485 ;
      RECT 0.09 1.695 0.505 2.21 ;
      RECT 0.09 1.695 1.8 1.865 ;
      RECT 1.47 1.415 1.8 1.865 ;
      RECT 0.09 0.685 0.26 2.21 ;
      RECT 0.09 0.685 0.355 1.015 ;
  END
END scs130lp_nand2b_2

MACRO scs130lp_nand2b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2b_4 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.365 0.495 1.76 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.25 1.425 5.18 1.76 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.016 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.295 1.93 4.515 3.075 ;
        RECT 2.365 1.93 4.515 2.1 ;
        RECT 3.36 1.93 3.69 3.075 ;
        RECT 2.365 1.93 3.69 2.12 ;
        RECT 1.435 1.765 3.08 1.935 ;
        RECT 2.62 1.44 3.08 2.12 ;
        RECT 2.62 0.605 2.805 2.12 ;
        RECT 2.365 1.765 2.665 3.075 ;
        RECT 1.475 1.085 2.805 1.255 ;
        RECT 2.475 0.605 2.805 1.255 ;
        RECT 1.475 0.605 1.805 1.255 ;
        RECT 1.435 1.765 1.695 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.195 -0.085 4.525 0.905 ;
        RECT 3.335 -0.085 3.665 0.915 ;
        RECT 0.525 -0.085 0.855 0.855 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.685 1.93 5.015 3.415 ;
        RECT 3.86 2.27 4.125 3.415 ;
        RECT 2.835 2.29 3.165 3.415 ;
        RECT 1.865 2.105 2.195 3.415 ;
        RECT 0.525 2.27 1.265 3.415 ;
        RECT 1.005 1.8 1.265 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.975 1.085 4.955 1.255 ;
      RECT 4.695 0.305 4.955 1.255 ;
      RECT 1.045 0.255 1.305 1.185 ;
      RECT 3.835 1.075 4.955 1.255 ;
      RECT 2.975 0.255 3.165 1.255 ;
      RECT 3.835 0.285 4.025 1.255 ;
      RECT 1.975 0.255 2.305 0.915 ;
      RECT 1.045 0.255 3.165 0.425 ;
      RECT 0.095 1.93 0.355 3.075 ;
      RECT 0.095 1.93 0.835 2.1 ;
      RECT 0.665 1.025 0.835 2.1 ;
      RECT 0.665 1.425 2.45 1.595 ;
      RECT 0.095 1.025 0.835 1.195 ;
      RECT 0.095 0.255 0.345 1.195 ;
  END
END scs130lp_nand2b_4

MACRO scs130lp_nand2b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2b_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.485 1.225 0.835 1.895 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.225 1.385 1.895 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3997 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.135 0.265 2.305 2.15 ;
        RECT 1.565 1.92 2.305 2.15 ;
        RECT 1.75 0.265 2.305 0.695 ;
        RECT 1.32 2.075 1.735 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.93 -0.085 1.26 0.695 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.915 2.33 2.245 3.415 ;
        RECT 0.79 2.075 1.12 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.135 2.075 0.59 3.065 ;
      RECT 0.135 0.265 0.305 3.065 ;
      RECT 1.625 0.875 1.955 1.545 ;
      RECT 0.135 0.875 1.955 1.045 ;
      RECT 0.135 0.265 0.47 1.045 ;
  END
END scs130lp_nand2b_lp

MACRO scs130lp_nand2b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand2b_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.62 0.47 0.805 2.12 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.8 1.33 1.47 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.335 2.48 2.245 2.65 ;
        RECT 2.075 0.44 2.245 2.65 ;
        RECT 1.745 0.44 2.245 0.65 ;
        RECT 1.335 2.48 1.525 2.97 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.985 -0.085 1.195 0.58 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.705 2.83 2.035 3.415 ;
        RECT 0.905 2.77 1.115 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.475 2.3 0.685 2.97 ;
      RECT 0.25 2.3 1.155 2.47 ;
      RECT 1.54 1.79 1.87 2.3 ;
      RECT 0.985 2.13 1.87 2.3 ;
      RECT 0.25 0.38 0.44 2.47 ;
  END
END scs130lp_nand2b_m

MACRO scs130lp_nand3_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3_0 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.095 0.84 1.475 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.57 0.78 0.925 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.355 2.12 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4601 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.44 1.92 1.835 2.97 ;
        RECT 1.645 0.28 1.835 2.97 ;
        RECT 1.34 0.28 1.835 0.61 ;
        RECT 0.585 1.92 1.835 2.12 ;
        RECT 0.585 1.92 0.84 2.97 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.13 -0.085 0.46 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.01 2.29 1.27 3.415 ;
        RECT 0.12 2.29 0.415 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand3_0

MACRO scs130lp_nand3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.51 0.47 1.765 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 0.47 1.34 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.855 1.75 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1151 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.665 1.92 2.315 3.075 ;
        RECT 1.935 0.36 2.315 3.075 ;
        RECT 0.635 1.92 2.315 2.12 ;
        RECT 0.635 1.92 0.995 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.25 -0.085 0.58 1.03 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.165 2.29 1.495 3.415 ;
        RECT 0.215 1.92 0.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand3_1

MACRO scs130lp_nand3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.505 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.49 1.425 3.05 1.645 ;
        RECT 1.105 1.92 2.745 2.12 ;
        RECT 2.49 1.425 2.745 2.12 ;
        RECT 1.105 1.425 1.6 2.12 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.81 1.425 2.32 1.75 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.455 2.29 2.745 3.075 ;
        RECT 1.555 2.29 2.745 2.49 ;
        RECT 1.555 2.29 1.785 3.075 ;
        RECT 0.675 2.29 2.745 2.46 ;
        RECT 0.675 0.595 0.935 2.46 ;
        RECT 0.675 0.595 0.885 3.075 ;
        RECT 0.605 0.595 0.935 1.07 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.985 -0.085 2.315 0.575 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.915 1.815 3.175 3.415 ;
        RECT 1.955 2.66 2.285 3.415 ;
        RECT 1.055 2.63 1.385 3.415 ;
        RECT 0.175 1.92 0.505 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.105 1.085 3.245 1.255 ;
      RECT 2.985 0.305 3.245 1.255 ;
      RECT 1.105 0.255 1.315 1.255 ;
      RECT 0.175 0.255 0.435 1.04 ;
      RECT 0.175 0.255 1.315 0.425 ;
      RECT 1.485 0.745 2.815 0.915 ;
      RECT 2.485 0.285 2.815 0.915 ;
      RECT 1.485 0.285 1.815 0.915 ;
  END
END scs130lp_nand3_2

MACRO scs130lp_nand3_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.395 1.31 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.2 1.425 5.54 1.705 ;
        RECT 2.795 1.92 5.43 2.12 ;
        RECT 5.2 1.425 5.43 2.12 ;
        RECT 2.795 1.425 3.18 2.12 ;
        RECT 2.17 1.425 3.18 1.605 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.39 1.425 4.93 1.75 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.975 2.29 5.165 3.075 ;
        RECT 2.365 2.29 5.165 2.46 ;
        RECT 4.105 2.29 4.305 3.075 ;
        RECT 3.225 2.29 3.415 3.075 ;
        RECT 2.365 1.775 2.625 2.46 ;
        RECT 2.365 1.775 2.545 3.075 ;
        RECT 1.495 1.775 2.625 1.945 ;
        RECT 1.495 1.425 2 1.945 ;
        RECT 1.495 0.595 1.71 1.945 ;
        RECT 1.505 0.595 1.695 3.075 ;
        RECT 0.645 1.92 1.695 2.1 ;
        RECT 0.595 1.055 1.71 1.225 ;
        RECT 1.485 0.595 1.71 1.225 ;
        RECT 0.645 1.92 0.835 3.075 ;
        RECT 0.595 0.595 0.815 1.225 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.475 -0.085 4.805 0.575 ;
        RECT 3.675 -0.085 3.945 0.575 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.335 2.29 5.665 3.415 ;
        RECT 4.475 2.63 4.805 3.415 ;
        RECT 3.585 2.63 3.915 3.415 ;
        RECT 2.725 2.63 3.055 3.415 ;
        RECT 1.865 2.115 2.195 3.415 ;
        RECT 1.005 2.27 1.335 3.415 ;
        RECT 0.145 1.92 0.475 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.88 1.085 5.665 1.255 ;
      RECT 5.405 0.265 5.665 1.255 ;
      RECT 0.125 0.255 0.425 1.145 ;
      RECT 2.775 0.645 3.005 1.255 ;
      RECT 1.88 0.255 2.105 1.255 ;
      RECT 0.985 0.255 1.315 0.885 ;
      RECT 0.125 0.255 2.105 0.425 ;
      RECT 3.175 0.745 5.235 0.915 ;
      RECT 4.93 0.7 5.235 0.915 ;
      RECT 2.275 0.255 2.605 0.915 ;
      RECT 4.065 0.7 4.355 0.915 ;
      RECT 3.175 0.255 3.505 0.915 ;
      RECT 2.275 0.255 3.505 0.425 ;
  END
END scs130lp_nand3_4

MACRO scs130lp_nand3_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.855 1.915 1.525 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 0.44 1.345 1.435 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.855 0.835 1.525 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6847 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.81 1.705 2.265 3.065 ;
        RECT 2.095 0.505 2.265 3.065 ;
        RECT 1.71 0.505 2.265 0.675 ;
        RECT 1.71 0.265 2.04 0.675 ;
        RECT 0.605 1.705 2.265 1.875 ;
        RECT 0.605 1.705 1.08 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.32 -0.085 0.65 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.28 2.055 1.61 3.415 ;
        RECT 0.175 2.025 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand3_lp

MACRO scs130lp_nand3_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.84 1.465 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 0.925 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.12 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3402 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.47 1.95 1.815 2.74 ;
        RECT 1.645 0.405 1.815 2.74 ;
        RECT 1.34 0.405 1.815 0.615 ;
        RECT 0.61 1.95 1.815 2.12 ;
        RECT 0.61 1.95 0.82 2.74 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.13 -0.085 0.46 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.04 2.3 1.25 3.415 ;
        RECT 0.18 2.3 0.39 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand3_m

MACRO scs130lp_nand3b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3b_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.505 1.425 0.875 1.75 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.425 1.915 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.425 1.375 1.75 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9093 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.31 1.92 2.795 3.075 ;
        RECT 2.545 0.275 2.795 3.075 ;
        RECT 2.205 0.275 2.795 0.915 ;
        RECT 1.35 1.92 2.795 2.09 ;
        RECT 1.35 1.92 1.635 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.82 -0.085 1.19 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.805 2.26 2.135 3.415 ;
        RECT 0.88 1.92 1.18 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.155 1.92 0.71 2.21 ;
      RECT 0.155 0.765 0.325 2.21 ;
      RECT 2.125 1.085 2.375 1.515 ;
      RECT 0.155 1.085 2.375 1.255 ;
      RECT 0.155 0.765 0.65 1.255 ;
  END
END scs130lp_nand3b_1

MACRO scs130lp_nand3b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3b_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.43 1.345 0.83 1.75 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.735 3.33 1.905 ;
        RECT 2.52 1.345 3.33 1.905 ;
        RECT 1.53 1.345 1.72 1.905 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.19 2.075 3.79 2.245 ;
        RECT 3.54 1.345 3.79 2.245 ;
        RECT 1.19 1.345 1.36 2.245 ;
        RECT 1 1.345 1.36 1.75 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4532 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.225 2.415 4.235 2.585 ;
        RECT 3.96 1.005 4.235 2.585 ;
        RECT 2.24 1.005 4.235 1.175 ;
        RECT 3.235 2.415 3.565 3.075 ;
        RECT 2.245 2.415 2.575 3.075 ;
        RECT 2.24 0.935 2.57 1.175 ;
        RECT 1.225 2.415 1.555 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.665 -0.085 3.995 0.835 ;
        RECT 0.775 -0.085 1.105 0.835 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.735 2.755 3.995 3.415 ;
        RECT 2.745 2.755 3.065 3.415 ;
        RECT 1.735 2.755 2.065 3.415 ;
        RECT 0.735 1.92 1.02 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.265 0.255 3.495 0.835 ;
      RECT 1.275 0.255 1.535 0.835 ;
      RECT 1.275 0.255 3.495 0.425 ;
      RECT 2.765 0.595 3.095 0.835 ;
      RECT 1.705 0.595 2.035 0.835 ;
      RECT 1.705 0.595 3.095 0.765 ;
      RECT 0.09 1.92 0.565 2.2 ;
      RECT 0.09 0.825 0.26 2.2 ;
      RECT 1.89 1.345 2.35 1.565 ;
      RECT 1.89 1.005 2.06 1.565 ;
      RECT 0.09 1.005 2.06 1.175 ;
      RECT 0.09 0.825 0.565 1.175 ;
  END
END scs130lp_nand3b_2

MACRO scs130lp_nand3b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3b_4 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 1.21 0.805 1.75 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.405 4.735 1.76 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.95 1.405 7.045 1.76 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 6 1.93 6.19 3.075 ;
        RECT 2.265 1.93 6.19 2.1 ;
        RECT 5.035 1.93 5.33 3.075 ;
        RECT 4.05 1.93 4.365 3.075 ;
        RECT 3.145 1.93 3.38 3.075 ;
        RECT 1.355 1.69 3.205 1.945 ;
        RECT 2.265 1.93 3.38 2.49 ;
        RECT 2.92 1.21 3.205 2.49 ;
        RECT 2.92 0.975 3.09 2.49 ;
        RECT 1.515 0.975 3.09 1.145 ;
        RECT 2.445 0.595 2.635 1.145 ;
        RECT 2.265 1.69 2.455 3.075 ;
        RECT 1.515 0.595 1.775 1.145 ;
        RECT 1.355 1.69 1.595 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 6.8 -0.085 7.095 1.095 ;
        RECT 5.905 -0.085 6.235 0.895 ;
        RECT 5.045 -0.085 5.375 0.885 ;
        RECT 0.565 -0.085 0.895 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.36 1.93 6.69 3.415 ;
        RECT 5.5 2.27 5.83 3.415 ;
        RECT 4.535 2.27 4.865 3.415 ;
        RECT 3.55 2.27 3.88 3.415 ;
        RECT 2.625 2.66 2.955 3.415 ;
        RECT 1.765 2.115 2.095 3.415 ;
        RECT 0.91 1.885 1.185 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.375 1.065 6.63 1.235 ;
      RECT 6.405 0.255 6.63 1.235 ;
      RECT 3.33 1.065 6.63 1.085 ;
      RECT 3.305 0.615 3.495 1.065 ;
      RECT 5.545 0.255 5.735 1.235 ;
      RECT 3.305 0.955 4.355 1.065 ;
      RECT 4.165 0.615 4.355 1.235 ;
      RECT 4.525 0.255 4.855 0.895 ;
      RECT 2.805 0.255 3.135 0.805 ;
      RECT 1.945 0.255 2.275 0.805 ;
      RECT 3.665 0.255 3.995 0.785 ;
      RECT 1.085 0.255 1.345 0.7 ;
      RECT 2.805 0.255 4.855 0.445 ;
      RECT 1.085 0.255 4.855 0.425 ;
      RECT 0.135 1.92 0.74 3.075 ;
      RECT 0.135 0.87 0.405 3.075 ;
      RECT 0.975 1.315 2.75 1.52 ;
      RECT 0.975 0.87 1.32 1.52 ;
      RECT 0.135 0.87 1.32 1.04 ;
      RECT 0.135 0.36 0.395 3.075 ;
  END
END scs130lp_nand3b_4

MACRO scs130lp_nand3b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3b_lp 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 0.265 2.755 0.67 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.99 1.55 1.32 1.92 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.55 2.275 1.88 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6847 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.255 2.1 1.585 3.065 ;
        RECT 0.1 0.44 1.315 1.02 ;
        RECT 0.1 2.1 1.585 2.27 ;
        RECT 0.1 2.085 0.525 3.065 ;
        RECT 0.1 0.44 0.27 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.535 -0.085 1.865 1.02 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.785 2.06 2.115 3.415 ;
        RECT 0.725 2.45 1.055 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.355 2.06 2.765 3.065 ;
      RECT 2.595 0.85 2.765 3.065 ;
      RECT 0.45 1.2 0.78 1.905 ;
      RECT 0.45 1.2 2.765 1.37 ;
      RECT 2.435 0.85 2.765 1.37 ;
  END
END scs130lp_nand3b_lp

MACRO scs130lp_nand3b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand3b_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.46 0.84 0.805 1.75 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 0.47 1.795 1.38 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 0.47 1.285 1.435 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3507 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 0.405 2.305 2.205 ;
        RECT 1.115 1.715 2.305 1.885 ;
        RECT 1.595 1.58 2.305 1.885 ;
        RECT 1.115 1.715 1.445 2.205 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.655 -0.085 0.825 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.625 2.065 1.795 3.415 ;
        RECT 0.765 2.375 1.795 2.545 ;
        RECT 0.87 2.375 1.04 3.415 ;
        RECT 0.765 2.065 0.935 2.545 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.255 2.715 0.7 3.045 ;
      RECT 0.255 2.125 0.585 3.045 ;
      RECT 0.11 0.405 0.28 2.335 ;
      RECT 0.11 0.405 0.475 0.615 ;
  END
END scs130lp_nand3b_m

MACRO scs130lp_nand4_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 0.78 2.425 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 0.375 1.855 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 0.375 1.35 1.75 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.715 2.12 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4781 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.945 1.92 2.795 2.13 ;
        RECT 2.595 0.28 2.795 2.13 ;
        RECT 2.28 0.28 2.795 0.61 ;
        RECT 1.805 1.92 2.065 2.96 ;
        RECT 0.945 1.92 1.205 2.96 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.34 -0.085 0.67 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.235 2.3 2.53 3.415 ;
        RECT 1.375 2.3 1.635 3.415 ;
        RECT 0.48 2.29 0.775 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand4_0

MACRO scs130lp_nand4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.47 2.295 1.515 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.555 0.47 1.765 1.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.47 1.285 1.515 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.805 1.435 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.134 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.755 2.685 1.925 ;
        RECT 2.475 0.425 2.685 1.925 ;
        RECT 1.8 1.755 2.245 2.825 ;
        RECT 0.635 1.755 2.245 2.12 ;
        RECT 0.635 1.755 0.91 2.825 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.27 -0.085 0.48 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.425 2.105 2.635 3.415 ;
        RECT 1.13 2.445 1.34 3.415 ;
        RECT 0.245 2.105 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand4_1

MACRO scs130lp_nand4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 1.425 4.715 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.425 3.335 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.165 2.33 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 1.345 0.845 1.64 ;
        RECT 0.625 1.345 0.805 2.12 ;
        RECT 0.555 1.345 0.805 1.67 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.5 1.075 4.215 1.245 ;
        RECT 3.885 0.595 4.215 1.245 ;
        RECT 3.815 1.92 4.075 3.075 ;
        RECT 1.835 1.92 4.075 2.09 ;
        RECT 2.74 1.92 3.035 3.075 ;
        RECT 0.975 1.755 2.835 1.925 ;
        RECT 2.015 1.605 2.835 2.09 ;
        RECT 2.5 1.075 2.835 2.09 ;
        RECT 1.835 1.755 2.015 3.075 ;
        RECT 0.975 1.755 1.165 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 0.735 -0.085 1.065 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.245 1.92 4.575 3.415 ;
        RECT 3.26 2.26 3.59 3.415 ;
        RECT 2.24 2.26 2.57 3.415 ;
        RECT 1.335 2.095 1.665 3.415 ;
        RECT 0.135 2.295 0.805 3.415 ;
        RECT 0.135 1.815 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.385 0.255 4.645 1.195 ;
      RECT 3.525 0.255 3.715 0.905 ;
      RECT 2.595 0.255 3.715 0.545 ;
      RECT 2.595 0.255 4.645 0.425 ;
      RECT 1.625 0.715 1.955 0.995 ;
      RECT 1.625 0.715 3.355 0.905 ;
      RECT 0.305 0.985 1.415 1.155 ;
      RECT 1.235 0.255 1.415 1.155 ;
      RECT 0.305 0.255 0.565 1.155 ;
      RECT 1.235 0.255 2.385 0.545 ;
  END
END scs130lp_nand4_2

MACRO scs130lp_nand4_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.22 1.425 8.005 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.98 1.425 6.01 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.425 3.45 1.75 ;
        RECT 2.2 1.38 3.45 1.75 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.425 1.765 1.75 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.2928 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.63 1.085 7.535 1.255 ;
        RECT 7.205 0.625 7.535 1.255 ;
        RECT 7.275 1.92 7.465 3.075 ;
        RECT 0.61 1.92 7.465 2.09 ;
        RECT 6.345 0.625 6.675 1.255 ;
        RECT 6.415 1.92 6.605 3.075 ;
        RECT 5.105 1.92 5.295 3.075 ;
        RECT 4.245 1.92 4.435 3.075 ;
        RECT 3.63 1.085 3.8 2.09 ;
        RECT 3.385 1.92 3.575 3.075 ;
        RECT 2.445 1.92 2.715 3.075 ;
        RECT 1.505 1.92 1.765 3.075 ;
        RECT 0.61 1.92 1.765 2.12 ;
        RECT 0.61 1.92 0.835 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 1.385 -0.085 1.715 0.915 ;
        RECT 0.525 -0.085 0.855 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.635 1.92 7.965 3.415 ;
        RECT 6.775 2.26 7.105 3.415 ;
        RECT 5.465 2.26 6.245 3.415 ;
        RECT 4.605 2.26 4.935 3.415 ;
        RECT 3.745 2.26 4.075 3.415 ;
        RECT 2.885 2.26 3.215 3.415 ;
        RECT 1.945 2.26 2.275 3.415 ;
        RECT 1.005 2.29 1.335 3.415 ;
        RECT 0.145 1.92 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 7.705 0.275 7.965 1.195 ;
      RECT 6.845 0.275 7.035 0.915 ;
      RECT 5.985 0.275 6.175 0.915 ;
      RECT 4.195 0.275 6.175 0.575 ;
      RECT 4.195 0.275 7.965 0.445 ;
      RECT 2.245 1.035 3.435 1.205 ;
      RECT 3.105 0.605 3.435 1.205 ;
      RECT 2.245 0.605 2.575 1.205 ;
      RECT 3.105 0.745 5.815 0.915 ;
      RECT 0.155 1.085 2.075 1.255 ;
      RECT 1.885 0.265 2.075 1.255 ;
      RECT 1.025 0.305 1.215 1.255 ;
      RECT 0.155 0.305 0.355 1.255 ;
      RECT 2.745 0.265 2.935 0.865 ;
      RECT 3.615 0.265 3.945 0.565 ;
      RECT 1.885 0.265 3.945 0.435 ;
  END
END scs130lp_nand4_4

MACRO scs130lp_nand4_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4_lp 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.33 1.11 2.755 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.47 0.44 1.8 1.435 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.9 0.44 1.29 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.825 0.55 1.495 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6797 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 0.265 2.755 0.675 ;
        RECT 1.735 1.675 2.15 3.065 ;
        RECT 1.98 0.265 2.15 3.065 ;
        RECT 0.665 1.675 2.15 1.845 ;
        RECT 0.665 1.675 0.995 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.205 -0.085 0.535 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.33 2.025 2.66 3.415 ;
        RECT 1.195 2.025 1.525 3.415 ;
        RECT 0.135 2.025 0.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand4_lp

MACRO scs130lp_nand4_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.84 2.425 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.47 1.855 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.47 1.285 1.75 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.715 2.12 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3549 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.97 1.95 2.775 2.12 ;
        RECT 2.605 0.33 2.775 2.12 ;
        RECT 2.38 0.33 2.775 0.66 ;
        RECT 1.83 1.95 2.245 2.96 ;
        RECT 0.97 1.95 1.18 2.96 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.34 -0.085 0.67 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.425 2.3 2.635 3.415 ;
        RECT 1.4 2.3 1.61 3.415 ;
        RECT 0.54 2.3 0.75 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nand4_m

MACRO scs130lp_nand4b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4b_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.52 1.185 0.89 1.515 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 0.37 2.39 1.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 0.37 1.825 1.515 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 1.185 1.36 1.515 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9282 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.33 2.035 3.275 2.205 ;
        RECT 3.02 0.255 3.275 2.205 ;
        RECT 2.725 0.255 3.275 1.095 ;
        RECT 2.295 2.035 2.555 3.075 ;
        RECT 1.33 2.035 1.615 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 0.795 -0.085 1.125 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.725 2.375 3.055 3.415 ;
        RECT 1.785 2.375 2.115 3.415 ;
        RECT 0.745 2.035 1.16 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.695 0.575 2.2 ;
      RECT 0.085 1.695 2.85 1.865 ;
      RECT 2.6 1.345 2.85 1.865 ;
      RECT 0.085 0.685 0.35 2.2 ;
      RECT 0.085 0.685 0.625 1.015 ;
  END
END scs130lp_nand4b_1

MACRO scs130lp_nand4b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4b_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.035 0.435 1.625 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.925 1.415 2.735 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.425 4.715 1.75 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.885 1.425 5.605 1.75 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.659 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.885 1.92 5.075 3.075 ;
        RECT 1.505 1.92 5.075 2.09 ;
        RECT 4.025 1.92 4.215 3.075 ;
        RECT 2.44 1.92 4.215 2.12 ;
        RECT 2.905 1.075 3.215 2.12 ;
        RECT 1.475 1.075 3.215 1.245 ;
        RECT 2.44 1.92 2.675 3.075 ;
        RECT 1.475 0.595 1.805 1.245 ;
        RECT 1.505 1.92 1.77 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.825 -0.085 5.155 0.915 ;
        RECT 0.525 -0.085 0.855 0.525 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.245 1.92 5.575 3.415 ;
        RECT 4.385 2.26 4.715 3.415 ;
        RECT 2.845 2.29 3.855 3.415 ;
        RECT 1.94 2.26 2.27 3.415 ;
        RECT 0.955 1.815 1.335 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.445 1.085 5.605 1.255 ;
      RECT 5.325 0.325 5.605 1.255 ;
      RECT 4.455 0.325 4.655 1.255 ;
      RECT 3.445 0.595 3.775 1.255 ;
      RECT 3.955 0.255 4.285 0.915 ;
      RECT 2.475 0.255 2.805 0.555 ;
      RECT 2.475 0.255 4.285 0.425 ;
      RECT 1.045 0.255 1.305 1.185 ;
      RECT 1.975 0.725 3.235 0.905 ;
      RECT 2.975 0.645 3.235 0.905 ;
      RECT 1.975 0.255 2.305 0.905 ;
      RECT 1.045 0.255 2.305 0.425 ;
      RECT 0.42 1.895 0.785 2.225 ;
      RECT 0.605 0.695 0.785 2.225 ;
      RECT 0.605 1.415 1.755 1.645 ;
      RECT 0.155 0.695 0.785 0.865 ;
      RECT 0.155 0.3 0.345 0.865 ;
  END
END scs130lp_nand4b_2

MACRO scs130lp_nand4b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4b_4 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.365 0.435 1.76 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.845 1.425 4.7 1.78 ;
        RECT 3.01 1.425 4.7 1.605 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.23 1.425 6.92 1.595 ;
        RECT 5.23 1.425 6.085 1.75 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.785 1.425 9.02 1.75 ;
        RECT 7.21 1.425 9.02 1.595 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.2928 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.215 1.93 8.405 3.075 ;
        RECT 7.355 1.93 8.405 2.1 ;
        RECT 7.355 1.765 7.535 3.075 ;
        RECT 6.255 1.765 7.615 1.935 ;
        RECT 6.125 1.92 6.425 3.075 ;
        RECT 3.185 1.95 6.425 2.12 ;
        RECT 4.88 1.92 6.425 2.12 ;
        RECT 5.265 1.92 5.455 3.075 ;
        RECT 4.88 1.075 5.05 2.12 ;
        RECT 1.51 1.075 5.05 1.255 ;
        RECT 4.065 1.95 4.255 3.075 ;
        RECT 3.185 1.775 3.67 2.12 ;
        RECT 3.185 1.775 3.395 3.075 ;
        RECT 1.345 1.775 3.67 1.945 ;
        RECT 2.405 0.595 2.595 1.255 ;
        RECT 2.285 1.775 2.515 3.075 ;
        RECT 1.51 0.595 1.735 1.255 ;
        RECT 1.345 1.775 1.615 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 8.195 -0.085 8.525 0.895 ;
        RECT 7.335 -0.085 7.665 0.905 ;
        RECT 0.525 -0.085 0.855 0.855 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 8.575 1.92 8.905 3.415 ;
        RECT 7.715 2.27 8.045 3.415 ;
        RECT 6.595 2.105 7.185 3.415 ;
        RECT 5.625 2.29 5.955 3.415 ;
        RECT 4.425 2.29 5.095 3.415 ;
        RECT 3.565 2.29 3.895 3.415 ;
        RECT 2.685 2.115 3.015 3.415 ;
        RECT 1.785 2.125 2.115 3.415 ;
        RECT 0.945 1.815 1.175 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.975 1.075 8.955 1.245 ;
      RECT 8.695 0.305 8.955 1.245 ;
      RECT 7.835 0.305 8.025 1.245 ;
      RECT 6.975 0.255 7.165 1.245 ;
      RECT 5.965 0.255 6.295 0.905 ;
      RECT 5.105 0.255 6.295 0.555 ;
      RECT 5.105 0.255 7.165 0.435 ;
      RECT 5.53 1.075 6.805 1.255 ;
      RECT 6.475 0.605 6.805 1.255 ;
      RECT 5.53 0.725 5.795 1.255 ;
      RECT 3.275 0.725 5.795 0.905 ;
      RECT 3.275 0.685 4.465 0.905 ;
      RECT 1.045 0.255 1.34 1.115 ;
      RECT 2.765 0.255 3.095 0.905 ;
      RECT 1.905 0.255 2.235 0.905 ;
      RECT 2.765 0.255 4.895 0.515 ;
      RECT 1.045 0.255 4.895 0.425 ;
      RECT 0.445 1.93 0.775 3.075 ;
      RECT 0.605 1.025 0.775 3.075 ;
      RECT 0.605 1.425 2.8 1.595 ;
      RECT 0.605 1.025 0.855 1.595 ;
      RECT 0.095 1.025 0.855 1.195 ;
      RECT 0.095 0.255 0.345 1.195 ;
  END
END scs130lp_nand4b_4

MACRO scs130lp_nand4b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4b_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.175 2.905 1.845 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.45 1.255 1.78 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.175 1.795 1.845 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.175 2.335 1.845 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6797 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.72 2.025 2.05 3.065 ;
        RECT 0.66 2.025 2.05 2.195 ;
        RECT 0.66 1.96 0.99 3.065 ;
        RECT 0.125 0.475 0.74 0.645 ;
        RECT 0.41 0.265 0.74 0.645 ;
        RECT 0.125 1.96 0.99 2.13 ;
        RECT 0.125 0.475 0.355 2.13 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.01 -0.085 2.34 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.25 2.025 2.58 3.415 ;
        RECT 1.19 2.375 1.52 3.415 ;
        RECT 0.13 2.31 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.8 2.025 3.255 3.065 ;
      RECT 3.085 0.825 3.255 3.065 ;
      RECT 0.535 0.825 0.865 1.155 ;
      RECT 0.535 0.825 3.255 0.995 ;
      RECT 2.88 0.265 3.21 0.995 ;
  END
END scs130lp_nand4b_lp

MACRO scs130lp_nand4b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4b_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.565 0.84 0.805 2.49 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.47 2.435 1.38 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.47 1.895 1.38 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 0.47 1.355 1.38 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.58 3.205 1.75 ;
        RECT 3.035 0.43 3.205 1.75 ;
        RECT 2.77 0.43 3.205 0.64 ;
        RECT 2.195 1.58 2.525 2.21 ;
        RECT 1.335 1.58 1.665 2.21 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 0.675 -0.085 0.845 0.57 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.705 2.07 2.895 3.415 ;
        RECT 1.845 2.07 2.015 3.415 ;
        RECT 0.985 2.07 1.155 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.165 2.72 0.805 3.05 ;
      RECT 0.165 0.43 0.385 3.05 ;
      RECT 0.165 0.43 0.495 0.64 ;
  END
END scs130lp_nand4b_m

MACRO scs130lp_nand4bb_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4bb_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.42 0.805 3.86 1.39 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.2 0.805 2.975 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 1.2 2.01 1.52 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 1.21 1.345 1.75 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9282 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.65 0.255 3.25 1.11 ;
        RECT 2.455 1.69 2.82 3.075 ;
        RECT 2.65 0.255 2.82 3.075 ;
        RECT 1.515 1.69 2.82 1.86 ;
        RECT 1.515 1.69 1.775 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.42 -0.085 3.695 0.635 ;
        RECT 1.015 -0.085 1.345 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.99 1.9 3.475 3.415 ;
        RECT 1.95 2.03 2.28 3.415 ;
        RECT 0.975 1.92 1.345 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.645 1.56 3.915 2.215 ;
      RECT 2.99 1.56 4.21 1.73 ;
      RECT 4.03 0.305 4.21 1.73 ;
      RECT 2.99 1.345 3.25 1.73 ;
      RECT 3.865 0.305 4.21 0.635 ;
      RECT 0.205 0.82 0.465 2.21 ;
      RECT 2.22 0.82 2.48 1.52 ;
      RECT 0.205 0.82 2.48 1.03 ;
  END
END scs130lp_nand4bb_1

MACRO scs130lp_nand4bb_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4bb_2 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 0.775 1.305 1.445 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 0.775 0.845 1.445 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.855 1.21 4.645 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.435 1.425 6.085 1.75 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.1252 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.905 1.92 5.475 3.075 ;
        RECT 4.905 1.605 5.265 3.075 ;
        RECT 3.42 1.605 5.265 1.775 ;
        RECT 4.045 1.605 4.235 3.075 ;
        RECT 2.325 1.74 4.235 1.92 ;
        RECT 3.42 1.035 3.685 1.92 ;
        RECT 2.21 1.035 3.685 1.205 ;
        RECT 3.185 1.74 3.375 3.075 ;
        RECT 2.325 1.74 2.515 3.075 ;
        RECT 2.21 0.595 2.435 1.205 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.355 -0.085 5.685 0.895 ;
        RECT 0.66 -0.085 0.99 0.555 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.645 1.92 5.975 3.415 ;
        RECT 4.405 1.945 4.735 3.415 ;
        RECT 3.545 2.09 3.875 3.415 ;
        RECT 2.685 2.105 3.015 3.415 ;
        RECT 1.825 2.685 2.155 3.415 ;
        RECT 0.56 1.965 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.995 1.065 6.115 1.235 ;
      RECT 5.855 0.255 6.115 1.235 ;
      RECT 4.995 0.255 5.185 1.235 ;
      RECT 4.065 0.255 5.185 0.465 ;
      RECT 1.815 0.255 2.015 1.095 ;
      RECT 2.605 0.255 2.935 0.825 ;
      RECT 2.605 0.255 3.875 0.465 ;
      RECT 1.815 0.255 3.875 0.425 ;
      RECT 0.965 2.345 2.155 2.515 ;
      RECT 1.985 1.375 2.155 2.515 ;
      RECT 0.965 1.625 1.135 2.515 ;
      RECT 0.085 1.625 0.39 2.24 ;
      RECT 0.085 1.625 1.135 1.795 ;
      RECT 0.085 0.275 0.295 2.24 ;
      RECT 1.985 1.375 3.25 1.57 ;
      RECT 0.085 0.275 0.49 0.605 ;
      RECT 1.305 1.845 1.815 2.175 ;
      RECT 1.475 1.325 1.815 2.175 ;
      RECT 1.475 0.275 1.645 2.175 ;
      RECT 1.16 0.275 1.645 0.605 ;
      RECT 3.115 0.635 4.825 0.865 ;
  END
END scs130lp_nand4bb_2

MACRO scs130lp_nand4bb_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4bb_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.445 1.21 0.865 1.75 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.21 1.285 1.75 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.27 1.2 8.005 1.515 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.21 1.2 9.925 1.515 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.2928 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.265 1.685 9.485 3.075 ;
        RECT 2.345 1.775 9.485 1.945 ;
        RECT 6.255 1.685 9.485 1.945 ;
        RECT 8.405 1.685 8.595 3.075 ;
        RECT 7.545 1.685 7.735 3.075 ;
        RECT 6.645 1.685 6.875 3.075 ;
        RECT 4.925 1.775 6.085 2.16 ;
        RECT 4.925 1.775 5.115 3.075 ;
        RECT 3.995 1.775 6.085 2.12 ;
        RECT 3.995 1.775 4.255 3.075 ;
        RECT 3.52 0.955 3.69 1.945 ;
        RECT 2.145 0.955 3.69 1.215 ;
        RECT 3.205 1.775 3.425 3.075 ;
        RECT 2.345 1.775 2.535 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.225 -0.085 9.555 0.69 ;
        RECT 8.365 -0.085 8.695 0.69 ;
        RECT 0.63 -0.085 0.96 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.655 1.815 9.955 3.415 ;
        RECT 8.765 2.115 9.095 3.415 ;
        RECT 7.905 2.115 8.235 3.415 ;
        RECT 7.045 2.115 7.375 3.415 ;
        RECT 5.285 2.33 6.475 3.415 ;
        RECT 6.255 2.125 6.475 3.415 ;
        RECT 4.425 2.29 4.755 3.415 ;
        RECT 3.595 2.115 3.825 3.415 ;
        RECT 2.705 2.115 3.035 3.415 ;
        RECT 1.845 2.68 2.175 3.415 ;
        RECT 0.63 2.68 0.96 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.28 0.86 9.925 1.03 ;
      RECT 9.725 0.255 9.925 1.03 ;
      RECT 8.865 0.255 9.045 1.03 ;
      RECT 7.995 0.255 8.195 1.03 ;
      RECT 6.28 0.7 7.345 1.03 ;
      RECT 4.245 1.055 6.1 1.245 ;
      RECT 5.93 0.31 6.1 1.245 ;
      RECT 5.115 0.96 6.1 1.245 ;
      RECT 4.245 0.885 4.445 1.245 ;
      RECT 5.115 0.86 5.305 1.245 ;
      RECT 7.515 0.31 7.775 0.69 ;
      RECT 5.93 0.31 7.775 0.52 ;
      RECT 1.06 1.92 1.68 2.17 ;
      RECT 1.5 0.615 1.68 2.17 ;
      RECT 3.87 1.415 5.9 1.605 ;
      RECT 3.87 0.615 4.04 1.605 ;
      RECT 1.13 0.325 1.33 1.04 ;
      RECT 1.13 0.615 4.04 0.785 ;
      RECT 4.615 0.255 4.945 0.885 ;
      RECT 5.475 0.255 5.76 0.79 ;
      RECT 1.6 0.255 4.945 0.445 ;
      RECT 1.6 0.255 5.76 0.425 ;
      RECT 0.085 1.93 0.45 2.94 ;
      RECT 0.085 2.34 2.02 2.51 ;
      RECT 1.85 1.385 2.02 2.51 ;
      RECT 0.085 0.325 0.275 2.94 ;
      RECT 1.85 1.385 3.34 1.605 ;
      RECT 0.085 0.325 0.46 1.04 ;
  END
END scs130lp_nand4bb_4

MACRO scs130lp_nand4bb_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4bb_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 0.855 0.835 1.525 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.765 3.72 1.085 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.49 1.615 2.82 2.15 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.615 3.36 2.15 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6797 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.725 2.33 3.055 3.065 ;
        RECT 1.355 2.33 3.055 2.52 ;
        RECT 2.045 1.94 2.275 2.52 ;
        RECT 1.6 1.94 2.275 2.11 ;
        RECT 1.465 0.265 1.795 0.675 ;
        RECT 1.6 0.265 1.77 2.11 ;
        RECT 1.355 2.29 1.685 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.035 -0.085 3.365 0.585 ;
        RECT 0.905 -0.085 1.235 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.255 2.33 3.585 3.415 ;
        RECT 1.885 2.7 2.215 3.415 ;
        RECT 0.825 2.075 1.155 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.825 1.265 4.205 3.065 ;
      RECT 4.035 0.295 4.205 3.065 ;
      RECT 1.95 1.09 2.28 1.76 ;
      RECT 1.95 1.265 4.205 1.435 ;
      RECT 3.875 0.295 4.205 0.585 ;
      RECT 0.115 1.725 0.625 3.065 ;
      RECT 0.115 1.725 1.42 1.895 ;
      RECT 1.09 1.225 1.42 1.895 ;
      RECT 0.115 0.265 0.285 3.065 ;
      RECT 0.115 0.265 0.445 0.675 ;
  END
END scs130lp_nand4bb_lp

MACRO scs130lp_nand4bb_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nand4bb_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 0.79 3.305 1.38 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.445 1.21 0.805 1.75 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 0.42 1.765 1.615 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.285 1.285 1.615 ;
        RECT 1.115 0.42 1.285 1.615 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3777 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.045 2.855 1.215 ;
        RECT 2.645 0.885 2.855 1.215 ;
        RECT 2.075 1.045 2.36 2.54 ;
        RECT 1.27 1.815 2.36 1.985 ;
        RECT 1.27 1.815 1.48 2.365 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.975 -0.085 3.305 0.485 ;
        RECT 0.605 -0.085 0.935 1.005 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.54 2.225 2.87 3.415 ;
        RECT 1.72 2.165 1.89 3.415 ;
        RECT 0.91 2.395 1.1 3.415 ;
        RECT 0.745 2.165 0.955 2.605 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.205 1.56 3.535 2.305 ;
      RECT 2.54 1.56 3.675 1.89 ;
      RECT 3.485 0.325 3.675 1.89 ;
      RECT 0.22 2.775 0.74 3.075 ;
      RECT 0.22 2.185 0.55 3.075 ;
      RECT 0.095 0.82 0.265 2.395 ;
      RECT 0.095 0.82 0.425 1.03 ;
  END
END scs130lp_nand4bb_m

MACRO scs130lp_nor2_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_0 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.455 2.225 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 0.84 1.355 2.225 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2872 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 2.395 1.295 3.075 ;
        RECT 0.625 0.385 0.885 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 1.055 -0.085 1.335 0.67 ;
        RECT 0.145 -0.085 0.455 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.145 2.395 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor2_0

MACRO scs130lp_nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_1 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.435 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.21 1.355 1.75 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5691 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.92 1.275 3.075 ;
        RECT 0.625 0.325 0.815 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 0.985 -0.085 1.315 1.04 ;
        RECT 0.125 -0.085 0.455 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.125 1.92 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor2_1

MACRO scs130lp_nor2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.43 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 1.425 1.525 1.75 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8232 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.695 1.075 1.875 2.1 ;
        RECT 1.46 0.255 1.765 1.255 ;
        RECT 1.38 1.92 1.72 2.735 ;
        RECT 0.61 1.085 1.875 1.255 ;
        RECT 0.61 0.255 0.79 1.255 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.935 -0.085 2.185 0.905 ;
        RECT 0.96 -0.085 1.29 0.905 ;
        RECT 0.1 -0.085 0.43 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.53 2.26 0.86 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.03 2.905 2.295 3.075 ;
      RECT 2.045 1.82 2.295 3.075 ;
      RECT 0.1 1.92 0.36 3.075 ;
      RECT 1.03 1.92 1.21 3.075 ;
      RECT 0.1 1.92 1.21 2.09 ;
  END
END scs130lp_nor2_2

MACRO scs130lp_nor2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_4 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 1.21 1.525 1.56 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.425 4.165 1.76 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.375 1.95 3.635 2.735 ;
        RECT 2.51 1.085 3.625 1.255 ;
        RECT 3.405 0.265 3.625 1.255 ;
        RECT 2.505 1.95 3.635 2.12 ;
        RECT 2.505 1.95 2.78 2.735 ;
        RECT 2.505 1.325 2.735 2.735 ;
        RECT 2.51 0.265 2.735 2.735 ;
        RECT 1.695 1.325 2.735 1.56 ;
        RECT 1.695 0.265 1.91 1.56 ;
        RECT 0.825 0.87 1.91 1.04 ;
        RECT 1.685 0.265 1.91 1.04 ;
        RECT 0.825 0.265 1.015 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.795 -0.085 4.095 1.14 ;
        RECT 2.905 -0.085 3.235 0.915 ;
        RECT 2.08 -0.085 2.34 1.155 ;
        RECT 1.185 -0.085 1.515 0.7 ;
        RECT 0.325 -0.085 0.655 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 1.615 2.095 1.945 3.415 ;
        RECT 0.755 2.095 1.085 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.115 2.905 4.095 3.075 ;
      RECT 3.805 1.93 4.095 3.075 ;
      RECT 1.255 1.73 1.445 3.075 ;
      RECT 0.325 1.73 0.585 3.075 ;
      RECT 2.95 2.29 3.205 3.075 ;
      RECT 2.115 1.73 2.335 3.075 ;
      RECT 0.325 1.73 2.335 1.925 ;
  END
END scs130lp_nor2_4

MACRO scs130lp_nor2_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_8 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.5 1.415 2.245 1.77 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.415 1.425 7.1 1.75 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.2928 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.065 1.92 7.595 2.09 ;
        RECT 7.425 1.085 7.595 2.09 ;
        RECT 4.995 1.085 7.595 1.255 ;
        RECT 6.645 1.92 6.975 2.725 ;
        RECT 6.715 0.305 6.905 1.255 ;
        RECT 5.785 1.92 6.115 2.725 ;
        RECT 5.855 0.305 6.045 1.255 ;
        RECT 4.925 1.92 5.255 2.735 ;
        RECT 4.065 1.36 5.245 2.09 ;
        RECT 4.995 1.085 5.245 2.735 ;
        RECT 4.995 0.305 5.185 2.735 ;
        RECT 4.065 1.36 4.395 2.735 ;
        RECT 2.425 1.21 4.325 1.485 ;
        RECT 4.135 0.305 4.325 2.735 ;
        RECT 3.275 0.305 3.465 1.485 ;
        RECT 0.68 1.075 2.605 1.245 ;
        RECT 2.415 0.305 2.605 1.245 ;
        RECT 1.555 0.315 1.745 1.245 ;
        RECT 0.68 0.315 0.885 1.245 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.075 -0.085 7.405 0.915 ;
        RECT 6.215 -0.085 6.545 0.915 ;
        RECT 5.355 -0.085 5.685 0.915 ;
        RECT 4.495 -0.085 4.825 1.19 ;
        RECT 3.635 -0.085 3.965 1.04 ;
        RECT 2.775 -0.085 3.105 1.04 ;
        RECT 1.915 -0.085 2.245 0.905 ;
        RECT 1.055 -0.085 1.385 0.905 ;
        RECT 0.185 -0.085 0.51 1.185 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 3.205 2.095 3.535 3.415 ;
        RECT 2.345 2.28 2.675 3.415 ;
        RECT 1.485 2.28 1.815 3.415 ;
        RECT 0.625 2.28 0.955 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.705 2.905 7.405 3.075 ;
      RECT 7.145 2.26 7.405 3.075 ;
      RECT 2.845 1.7 3.035 3.075 ;
      RECT 1.985 1.94 2.175 3.075 ;
      RECT 1.125 1.94 1.315 3.075 ;
      RECT 0.185 1.94 0.455 3.075 ;
      RECT 5.425 2.895 7.405 3.075 ;
      RECT 4.565 2.26 4.755 3.075 ;
      RECT 3.705 1.7 3.895 3.075 ;
      RECT 6.285 2.26 6.475 3.075 ;
      RECT 5.425 2.26 5.615 3.075 ;
      RECT 0.185 1.94 3.035 2.11 ;
      RECT 2.83 1.7 3.035 2.11 ;
      RECT 2.83 1.7 3.895 1.925 ;
  END
END scs130lp_nor2_8

MACRO scs130lp_nor2_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 2.15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.18 2.275 2.89 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2373 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 0.44 1.345 2.89 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.835 -0.085 2.165 1 ;
        RECT 0.195 -0.085 0.525 1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.195 2.43 0.525 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor2_lp

MACRO scs130lp_nor2_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_lp2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.18 2.275 2.89 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3826 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 0.44 1.395 2.89 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.835 -0.085 2.165 1 ;
        RECT 0.195 -0.085 0.525 1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.115 1.98 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor2_lp2

MACRO scs130lp_nor2_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2_m 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.455 2.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 0.84 1.285 2.12 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 2.395 1.235 2.845 ;
        RECT 0.635 0.33 0.885 2.86 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.44 0.085 ;
        RECT 1.065 -0.085 1.275 0.66 ;
        RECT 0.205 -0.085 0.415 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.44 3.415 ;
        RECT 0.205 2.405 0.415 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor2_m

MACRO scs130lp_nor2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2b_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.425 1.415 1.75 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.425 0.865 1.75 ;
    END
  END BN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8526 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.925 1.815 2.315 3.075 ;
        RECT 2.055 0.745 2.315 3.075 ;
        RECT 1.39 0.745 2.315 0.915 ;
        RECT 1.39 0.255 1.65 0.915 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.82 -0.085 2.15 0.575 ;
        RECT 0.795 -0.085 1.22 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.96 2.31 1.29 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.42 1.92 1.755 2.14 ;
      RECT 1.585 1.085 1.755 2.14 ;
      RECT 1.585 1.085 1.885 1.515 ;
      RECT 0.355 1.085 1.885 1.255 ;
      RECT 0.355 0.285 0.625 1.255 ;
  END
END scs130lp_nor2b_1

MACRO scs130lp_nor2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2b_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.075 2.815 1.515 ;
        RECT 1.055 1.075 2.815 1.245 ;
        RECT 1.055 1.075 1.775 1.435 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.6 1.185 0.885 1.515 ;
    END
  END BN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8232 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.82 2.025 3.275 2.195 ;
        RECT 2.985 0.735 3.275 2.195 ;
        RECT 1.435 0.735 3.275 0.905 ;
        RECT 2.365 0.255 2.555 0.905 ;
        RECT 1.82 2.025 2.15 2.715 ;
        RECT 1.435 0.255 1.695 0.905 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.725 -0.085 3.055 0.565 ;
        RECT 1.865 -0.085 2.195 0.565 ;
        RECT 0.62 -0.085 1.265 0.885 ;
        RECT 0.62 -0.085 0.895 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.68 2.365 3.01 3.415 ;
        RECT 0.865 2.025 1.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.42 2.895 2.51 3.075 ;
      RECT 2.32 2.365 2.51 3.075 ;
      RECT 1.42 2.025 1.65 3.075 ;
      RECT 0.16 1.685 0.695 2.21 ;
      RECT 0.16 1.685 2.275 1.855 ;
      RECT 1.945 1.415 2.275 1.855 ;
      RECT 0.16 0.7 0.43 2.21 ;
  END
END scs130lp_nor2b_2

MACRO scs130lp_nor2b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2b_4 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.965 1.695 4.305 1.865 ;
        RECT 4.045 1.345 4.305 1.865 ;
        RECT 2.065 1.425 3.205 1.865 ;
        RECT 0.965 1.425 1.295 1.865 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.345 0.435 1.76 ;
    END
  END BN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.63 2.035 4.7 2.205 ;
        RECT 4.475 1.005 4.7 2.205 ;
        RECT 3.84 1.005 4.7 1.175 ;
        RECT 3.84 0.745 4.03 1.175 ;
        RECT 3.85 0.255 4.03 1.175 ;
        RECT 1.2 0.745 4.03 0.915 ;
        RECT 3.41 2.035 3.62 2.715 ;
        RECT 2.92 0.255 3.25 0.915 ;
        RECT 2.06 0.255 2.39 0.915 ;
        RECT 1.63 2.035 1.96 2.255 ;
        RECT 1.2 0.255 1.53 0.915 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.21 -0.085 4.54 0.835 ;
        RECT 3.42 -0.085 3.68 0.575 ;
        RECT 2.56 -0.085 2.75 0.575 ;
        RECT 1.7 -0.085 1.89 0.575 ;
        RECT 0.69 -0.085 1.02 0.835 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.21 2.375 4.54 3.415 ;
        RECT 0.75 2.425 2.82 2.655 ;
        RECT 0.75 2.27 1.08 2.655 ;
        RECT 0.75 2.27 1.03 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.2 2.885 4.04 3.065 ;
      RECT 3.84 2.375 4.04 3.065 ;
      RECT 1.2 2.825 3.19 3.065 ;
      RECT 2.99 2.375 3.19 3.065 ;
      RECT 0.26 1.93 0.53 3.075 ;
      RECT 0.26 1.93 0.785 2.1 ;
      RECT 0.615 1.005 0.785 2.1 ;
      RECT 3.375 1.085 3.635 1.515 ;
      RECT 1.565 1.085 1.895 1.515 ;
      RECT 0.615 1.085 3.635 1.255 ;
      RECT 0.26 1.005 0.785 1.175 ;
      RECT 0.26 0.255 0.52 1.175 ;
  END
END scs130lp_nor2b_4

MACRO scs130lp_nor2b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2b_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 1.315 1.78 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.175 2.875 1.845 ;
    END
  END BN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 2.02 2.07 3.06 ;
        RECT 1.565 0.265 1.795 3.06 ;
        RECT 1.31 0.265 1.795 0.725 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.1 -0.085 2.43 0.645 ;
        RECT 0.52 -0.085 0.85 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.36 2.025 2.69 3.415 ;
        RECT 0.72 2.02 1.05 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.89 2.025 3.225 3.065 ;
      RECT 3.055 0.265 3.225 3.065 ;
      RECT 1.975 0.825 2.305 1.84 ;
      RECT 1.975 0.825 3.225 0.995 ;
      RECT 2.89 0.265 3.225 0.995 ;
  END
END scs130lp_nor2b_lp

MACRO scs130lp_nor2b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor2b_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.84 1.335 2.12 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.47 0.805 2.12 ;
    END
  END BN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.055 0.84 2.245 2.86 ;
        RECT 1.515 0.84 2.245 1.01 ;
        RECT 1.515 0.45 1.685 1.01 ;
        RECT 1.335 0.45 1.685 0.66 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.865 -0.085 2.055 0.66 ;
        RECT 0.985 -0.085 1.155 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.09 2.65 1.42 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.58 2.3 0.91 2.71 ;
      RECT 0.255 2.3 1.875 2.47 ;
      RECT 1.705 1.29 1.875 2.47 ;
      RECT 0.255 0.46 0.445 2.47 ;
  END
END scs130lp_nor2b_m

MACRO scs130lp_nor3_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3_0 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.405 2.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.21 0.925 2.86 ;
        RECT 0.575 1.21 0.925 2.215 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.095 1.21 1.465 2.2 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3985 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.37 2.395 1.835 3.065 ;
        RECT 1.635 0.365 1.835 3.065 ;
        RECT 0.575 0.84 1.835 1.04 ;
        RECT 1.48 0.365 1.835 1.04 ;
        RECT 0.575 0.79 0.81 1.04 ;
        RECT 0.62 0.365 0.81 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.98 -0.085 1.31 0.67 ;
        RECT 0.12 -0.085 0.45 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.16 2.405 0.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor3_0

MACRO scs130lp_nor3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3_1 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.455 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.345 1.01 1.68 ;
        RECT 0.625 1.345 0.905 2.925 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.21 1.835 1.675 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7917 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.425 1.845 1.835 3.075 ;
        RECT 0.595 0.87 1.755 1.04 ;
        RECT 1.475 0.255 1.755 1.04 ;
        RECT 1.18 1.845 1.835 2.165 ;
        RECT 1.18 0.87 1.35 2.165 ;
        RECT 0.595 0.255 0.805 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.975 -0.085 1.305 0.7 ;
        RECT 0.095 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.095 1.92 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor3_1

MACRO scs130lp_nor3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.185 1.16 1.515 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.67 1.605 3.745 1.785 ;
        RECT 2.94 1.285 3.745 1.785 ;
        RECT 1.67 1.345 1.87 1.785 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.04 1.21 2.76 1.435 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1172 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.33 0.84 2.98 1.04 ;
        RECT 2.755 0.255 2.98 1.04 ;
        RECT 1.33 1.965 2.505 2.295 ;
        RECT 1.845 0.255 2.085 1.04 ;
        RECT 1.33 0.84 1.5 2.295 ;
        RECT 0.965 0.84 2.98 1.015 ;
        RECT 0.965 0.255 1.175 1.015 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.15 -0.085 3.445 1.095 ;
        RECT 2.255 -0.085 2.585 0.67 ;
        RECT 1.345 -0.085 1.675 0.67 ;
        RECT 0.465 -0.085 0.795 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 0.58 2.815 1.245 3.415 ;
        RECT 0.58 2.025 0.82 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.485 1.955 3.745 3.075 ;
      RECT 1.415 2.465 1.605 3.075 ;
      RECT 0.14 1.685 0.41 3.075 ;
      RECT 0.99 2.465 2.845 2.645 ;
      RECT 2.675 1.955 2.845 2.645 ;
      RECT 0.99 1.685 1.16 2.645 ;
      RECT 2.675 1.955 3.745 2.125 ;
      RECT 0.14 1.685 1.16 1.855 ;
      RECT 1.775 2.815 3.315 3.075 ;
      RECT 3.015 2.295 3.315 3.075 ;
  END
END scs130lp_nor3_2

MACRO scs130lp_nor3_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 1.21 1.85 1.515 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.07 1.075 5.33 1.515 ;
        RECT 3.035 1.075 5.33 1.245 ;
        RECT 2.02 1.21 3.25 1.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.42 1.415 4.77 1.645 ;
        RECT 3.42 1.415 4.235 1.765 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.1168 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.5 0.725 5.67 1.985 ;
        RECT 4.405 1.815 5.67 1.985 ;
        RECT 2.325 0.725 5.67 0.895 ;
        RECT 4.835 0.255 5.165 0.895 ;
        RECT 3.545 1.935 4.735 2.155 ;
        RECT 3.975 0.255 4.305 0.895 ;
        RECT 3.115 0.255 3.445 0.895 ;
        RECT 0.575 0.87 2.865 1.04 ;
        RECT 2.325 0.255 2.545 1.04 ;
        RECT 1.465 0.255 1.655 1.04 ;
        RECT 0.575 0.255 0.795 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 5.335 -0.085 5.595 0.555 ;
        RECT 4.475 -0.085 4.665 0.555 ;
        RECT 3.615 -0.085 3.805 0.555 ;
        RECT 2.715 -0.085 2.945 0.555 ;
        RECT 1.825 -0.085 2.155 0.7 ;
        RECT 0.965 -0.085 1.295 0.7 ;
        RECT 0.105 -0.085 0.405 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 1.395 2.105 1.725 3.415 ;
        RECT 0.535 2.105 0.865 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.285 2.155 5.615 3.075 ;
      RECT 1.895 1.705 2.085 3.075 ;
      RECT 1.035 1.705 1.225 3.075 ;
      RECT 0.105 1.705 0.365 3.075 ;
      RECT 2.755 2.325 5.615 2.495 ;
      RECT 2.755 1.705 3.015 2.495 ;
      RECT 0.105 1.705 3.015 1.875 ;
      RECT 2.255 2.675 5.105 3.075 ;
      RECT 2.255 2.055 2.585 3.075 ;
  END
END scs130lp_nor3_4

MACRO scs130lp_nor3_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.005 3.235 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.18 2.275 2.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.175 1.385 1.845 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5223 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 0.265 2.32 0.725 ;
        RECT 0.41 0.825 2.16 0.995 ;
        RECT 1.99 0.265 2.16 0.995 ;
        RECT 0.93 2.025 1.26 3.065 ;
        RECT 0.125 2.025 1.26 2.89 ;
        RECT 0.125 1.18 0.835 2.89 ;
        RECT 0.41 0.825 0.835 2.89 ;
        RECT 0.41 0.265 0.74 2.89 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.78 -0.085 3.11 0.725 ;
        RECT 1.2 -0.085 1.53 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.52 2.025 2.85 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor3_lp

MACRO scs130lp_nor3_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.21 0.925 2.86 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.21 1.465 2.12 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3402 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.43 2.395 1.815 2.845 ;
        RECT 1.645 0.435 1.815 2.845 ;
        RECT 0.61 0.84 1.815 1.01 ;
        RECT 1.47 0.435 1.815 1.01 ;
        RECT 0.61 0.435 0.82 1.01 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.04 -0.085 1.25 0.635 ;
        RECT 0.18 -0.085 0.39 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 0.185 2.405 0.395 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor3_m

MACRO scs130lp_nor3b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3b_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 1.34 1.36 1.76 ;
        RECT 1.03 1.18 1.285 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.345 1.835 1.755 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.475 1.21 0.86 1.76 ;
    END
  END CN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.84 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.345 1.84 2.795 3.075 ;
        RECT 2.555 0.255 2.795 3.075 ;
        RECT 1.455 1 2.795 1.17 ;
        RECT 2.315 0.255 2.795 1.17 ;
        RECT 1.455 0.255 1.645 1.17 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.815 -0.085 2.145 0.83 ;
        RECT 0.8 -0.085 1.25 1.01 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 0.92 2.31 1.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.93 2.175 2.14 ;
      RECT 2.005 1.34 2.175 2.14 ;
      RECT 0.085 0.7 0.305 2.14 ;
      RECT 2.005 1.34 2.385 1.67 ;
      RECT 0.085 0.7 0.63 1.03 ;
  END
END scs130lp_nor3b_1

MACRO scs130lp_nor3b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3b_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.335 4.715 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.86 1.335 3.215 1.75 ;
        RECT 2.44 1.335 3.215 1.665 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.45 0.47 2.13 ;
    END
  END CN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1466 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.995 3.75 1.165 ;
        RECT 3.52 0.255 3.75 1.165 ;
        RECT 1.595 0.985 2.85 1.165 ;
        RECT 2.62 0.255 2.85 1.165 ;
        RECT 1.595 0.255 1.925 1.165 ;
        RECT 1.475 1.845 1.805 2.735 ;
        RECT 1.595 0.255 1.805 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.92 -0.085 4.21 1.095 ;
        RECT 3.02 -0.085 3.35 0.825 ;
        RECT 2.12 -0.085 2.45 0.815 ;
        RECT 0.525 -0.085 1.425 0.94 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.37 1.92 4.7 3.415 ;
        RECT 3.51 2.26 3.84 3.415 ;
        RECT 0.525 2.64 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.01 1.92 4.19 3.075 ;
      RECT 2.335 1.845 2.665 2.735 ;
      RECT 2.335 1.92 4.19 2.09 ;
      RECT 1.095 2.905 3.095 3.075 ;
      RECT 2.835 2.26 3.095 3.075 ;
      RECT 1.975 1.805 2.165 3.075 ;
      RECT 1.095 1.805 1.305 3.075 ;
      RECT 0.095 2.3 0.355 2.915 ;
      RECT 0.095 2.3 0.925 2.47 ;
      RECT 0.755 1.11 0.925 2.47 ;
      RECT 0.755 1.185 1.425 1.515 ;
      RECT 0.095 1.11 0.925 1.28 ;
      RECT 0.095 0.7 0.355 1.28 ;
  END
END scs130lp_nor3b_2

MACRO scs130lp_nor3b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3b_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 1.355 2.685 1.525 ;
        RECT 1.115 1.325 2.685 1.525 ;
        RECT 1.115 1.185 1.955 1.525 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.865 1.335 6.215 1.505 ;
        RECT 4.865 1.21 5.67 1.505 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.445 1.185 0.825 1.515 ;
    END
  END CN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.1168 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.33 1.675 6.635 1.855 ;
        RECT 6.385 0.985 6.635 1.855 ;
        RECT 5.84 0.985 6.635 1.155 ;
        RECT 4 0.87 6.04 1.04 ;
        RECT 5.85 0.255 6.04 1.155 ;
        RECT 4.925 0.255 5.18 1.04 ;
        RECT 3.33 1.675 4.4 2.145 ;
        RECT 2.21 0.985 4.26 1.155 ;
        RECT 4 0.255 4.255 1.155 ;
        RECT 3.14 0.255 3.33 1.155 ;
        RECT 1.305 0.845 2.47 1.015 ;
        RECT 2.24 0.255 2.47 1.155 ;
        RECT 1.305 0.255 1.57 1.015 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 6.21 -0.085 6.54 0.815 ;
        RECT 5.35 -0.085 5.68 0.7 ;
        RECT 4.425 -0.085 4.755 0.7 ;
        RECT 3.5 -0.085 3.83 0.815 ;
        RECT 2.64 -0.085 2.97 0.815 ;
        RECT 1.74 -0.085 2.07 0.675 ;
        RECT 0.805 -0.085 1.135 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 2.32 2.665 2.65 3.415 ;
        RECT 1.46 2.395 1.79 3.415 ;
        RECT 0.6 2.105 0.93 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.9 2.885 6.61 3.075 ;
      RECT 6.35 2.025 6.61 3.075 ;
      RECT 2.9 2.875 5.68 3.075 ;
      RECT 5.49 2.375 5.68 3.075 ;
      RECT 2.9 2.665 4.03 3.075 ;
      RECT 1.96 2.045 2.15 3.065 ;
      RECT 1.1 2.045 1.29 3.065 ;
      RECT 5.85 2.025 6.18 2.705 ;
      RECT 4.99 2.025 5.32 2.705 ;
      RECT 1.96 2.325 5.32 2.495 ;
      RECT 1.96 2.045 2.22 2.495 ;
      RECT 1.1 2.045 2.22 2.225 ;
      RECT 4.99 2.025 6.18 2.205 ;
      RECT 0.095 1.705 0.42 3.075 ;
      RECT 0.095 1.705 3.065 1.875 ;
      RECT 2.895 1.325 3.065 1.875 ;
      RECT 0.095 0.255 0.275 3.075 ;
      RECT 2.895 1.325 4.585 1.505 ;
      RECT 0.095 0.255 0.58 1.015 ;
  END
END scs130lp_nor3b_4

MACRO scs130lp_nor3b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3b_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.175 0.86 1.845 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.18 1.795 2.89 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.175 3.235 1.845 ;
    END
  END CN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5223 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 2.025 2.305 3.065 ;
        RECT 1.975 0.265 2.145 3.065 ;
        RECT 0.125 0.825 2.145 0.995 ;
        RECT 1.805 0.265 2.145 0.995 ;
        RECT 0.125 0.44 0.835 0.995 ;
        RECT 0.125 0.265 0.555 0.995 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.595 -0.085 2.925 0.645 ;
        RECT 1.015 -0.085 1.345 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.855 2.025 3.185 3.415 ;
        RECT 0.385 2.025 0.715 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.385 2.025 3.715 3.065 ;
      RECT 3.545 0.265 3.715 3.065 ;
      RECT 2.325 0.825 2.655 1.495 ;
      RECT 2.325 0.825 3.715 0.995 ;
      RECT 3.385 0.265 3.715 0.995 ;
  END
END scs130lp_nor3b_lp

MACRO scs130lp_nor3b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor3b_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.945 1.105 1.335 1.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.505 1.18 1.815 1.8 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.16 0.435 1.885 ;
    END
  END CN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3402 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 0.265 2.305 2.505 ;
        RECT 1.505 0.745 2.305 1.01 ;
        RECT 1.115 0.745 2.305 0.935 ;
        RECT 1.115 0.475 1.445 0.935 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.625 -0.085 1.835 0.575 ;
        RECT 0.745 -0.085 0.935 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 0.595 2.395 0.925 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.655 2.78 1.99 3.075 ;
      RECT 1.655 2.055 1.825 3.075 ;
      RECT 0.11 2.055 0.425 2.505 ;
      RECT 0.11 2.055 1.825 2.225 ;
      RECT 0.605 0.82 0.775 2.225 ;
      RECT 0.255 0.82 0.775 0.99 ;
      RECT 0.255 0.33 0.525 0.99 ;
  END
END scs130lp_nor3b_m

MACRO scs130lp_nor4_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.43 1.19 0.84 1.86 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 1.19 1.365 1.86 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.19 1.83 1.86 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 0.88 2.795 2.6 ;
        RECT 2.33 0.88 2.795 1.845 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4048 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 2.055 2.345 3.065 ;
        RECT 0.085 0.84 2.085 1.02 ;
        RECT 1.895 0.395 2.085 1.02 ;
        RECT 0.085 2.055 2.345 2.225 ;
        RECT 0.695 0.395 0.88 1.02 ;
        RECT 0.085 0.84 0.26 2.225 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.255 -0.085 2.585 0.71 ;
        RECT 1.05 -0.085 1.725 0.67 ;
        RECT 0.195 -0.085 0.525 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 0.415 2.405 0.745 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor4_0

MACRO scs130lp_nor4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.345 0.465 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.425 1.09 1.9 ;
        RECT 0.595 1.92 0.92 2.91 ;
        RECT 0.635 1.425 0.92 2.91 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.41 1.425 1.77 2.91 ;
        RECT 1.3 1.425 1.77 1.71 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.28 1.065 2.725 1.76 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8043 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.94 1.93 2.365 3.075 ;
        RECT 1.94 1.065 2.11 3.075 ;
        RECT 0.595 1.065 2.11 1.235 ;
        RECT 1.605 0.255 1.865 1.235 ;
        RECT 0.595 0.255 0.855 1.235 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.035 -0.085 2.365 0.895 ;
        RECT 1.065 -0.085 1.395 0.895 ;
        RECT 0.095 -0.085 0.425 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 0.095 1.92 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor4_1

MACRO scs130lp_nor4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.21 1.45 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.615 2.185 1.785 ;
        RECT 1.855 1.425 2.185 1.785 ;
        RECT 0.085 1.345 0.855 1.785 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.395 1.695 4.23 1.865 ;
        RECT 3.465 1.425 4.23 1.865 ;
        RECT 2.395 1.425 2.725 1.865 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.99 1.185 3.295 1.515 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.17 2.035 4.715 2.205 ;
        RECT 4.4 1.005 4.715 2.205 ;
        RECT 3.59 1.005 4.715 1.175 ;
        RECT 2.65 0.845 3.79 1.015 ;
        RECT 3.6 0.255 3.79 1.175 ;
        RECT 3.17 2.035 3.5 2.335 ;
        RECT 2.65 0.255 2.93 1.015 ;
        RECT 1.62 1.085 2.82 1.255 ;
        RECT 2.65 0.255 2.82 1.255 ;
        RECT 1.62 0.87 1.95 1.255 ;
        RECT 1.69 0.255 1.95 1.255 ;
        RECT 0.795 0.87 1.95 1.04 ;
        RECT 0.795 0.265 1.01 1.04 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.96 -0.085 4.29 0.835 ;
        RECT 3.1 -0.085 3.43 0.675 ;
        RECT 2.15 -0.085 2.48 0.915 ;
        RECT 1.19 -0.085 1.52 0.7 ;
        RECT 0.33 -0.085 0.625 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 1.19 2.635 1.52 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.085 2.905 4.36 3.075 ;
      RECT 4.1 2.375 4.36 3.075 ;
      RECT 0.33 1.955 0.625 3.075 ;
      RECT 2.085 2.035 2.53 3.075 ;
      RECT 0.33 1.955 2.24 2.125 ;
      RECT 2.74 2.505 3.93 2.735 ;
      RECT 2.74 2.035 3 2.735 ;
      RECT 1.69 2.295 1.915 3.075 ;
      RECT 0.795 2.295 1.02 3.075 ;
      RECT 0.795 2.295 1.915 2.465 ;
  END
END scs130lp_nor4_2

MACRO scs130lp_nor4_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.345 2.135 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.345 1.21 4.375 1.535 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.675 1.21 6.085 1.535 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.305 1.355 7.655 1.525 ;
        RECT 6.305 1.21 7.145 1.525 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.5 1.695 8.07 1.875 ;
        RECT 7.825 1.005 8.07 1.875 ;
        RECT 7.315 1.005 8.07 1.185 ;
        RECT 7.36 1.695 7.55 2.735 ;
        RECT 1.75 0.87 7.55 1.04 ;
        RECT 7.36 0.255 7.55 1.185 ;
        RECT 6.5 1.695 6.69 2.735 ;
        RECT 6.5 0.265 6.69 1.04 ;
        RECT 5.64 0.265 5.83 1.04 ;
        RECT 4.78 0.265 4.97 1.04 ;
        RECT 3.92 0.265 4.11 1.04 ;
        RECT 3.055 0.265 3.25 1.04 ;
        RECT 1.75 0.255 1.94 1.04 ;
        RECT 0.865 1.005 1.93 1.175 ;
        RECT 0.865 0.255 1.08 1.175 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.72 -0.085 8.05 0.835 ;
        RECT 6.86 -0.085 7.19 0.7 ;
        RECT 6 -0.085 6.33 0.7 ;
        RECT 5.14 -0.085 5.47 0.7 ;
        RECT 4.28 -0.085 4.61 0.7 ;
        RECT 3.42 -0.085 3.75 0.7 ;
        RECT 2.11 -0.085 2.885 0.7 ;
        RECT 1.25 -0.085 1.58 0.835 ;
        RECT 0.39 -0.085 0.695 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 1.61 2.26 1.94 3.415 ;
        RECT 0.75 2.26 1.08 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.28 2.905 8.05 3.075 ;
      RECT 7.72 2.055 8.05 3.075 ;
      RECT 6.86 2.055 7.19 3.075 ;
      RECT 6 2.055 6.33 3.075 ;
      RECT 5.14 2.055 5.47 3.075 ;
      RECT 4.28 2.055 4.61 3.075 ;
      RECT 5.64 1.705 5.82 2.735 ;
      RECT 4.78 1.705 4.97 2.735 ;
      RECT 3.4 1.705 3.615 2.725 ;
      RECT 2.515 1.705 2.73 2.725 ;
      RECT 2.515 1.705 5.82 1.875 ;
      RECT 2.11 2.895 4.09 3.065 ;
      RECT 3.785 2.055 4.09 3.065 ;
      RECT 1.25 1.92 1.44 3.065 ;
      RECT 0.32 1.92 0.58 3.065 ;
      RECT 2.9 2.055 3.23 3.065 ;
      RECT 2.11 1.92 2.345 3.065 ;
      RECT 0.32 1.92 2.345 2.09 ;
  END
END scs130lp_nor4_4

MACRO scs130lp_nor4_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.19 0.905 3.715 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.48 1.175 2.81 1.845 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.835 1.78 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.51 1.125 2.275 1.455 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5202 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 0.775 2.935 0.945 ;
        RECT 2.605 0.265 2.935 0.945 ;
        RECT 1.025 1.635 1.535 1.965 ;
        RECT 1.025 0.265 1.355 0.945 ;
        RECT 1.025 0.265 1.315 1.965 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.395 -0.085 3.725 0.725 ;
        RECT 1.815 -0.085 2.145 0.595 ;
        RECT 0.235 -0.085 0.565 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.315 2.025 3.645 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.645 2.895 2.625 3.065 ;
      RECT 2.295 2.025 2.625 3.065 ;
      RECT 0.645 2.495 0.975 3.065 ;
      RECT 0.115 2.025 0.445 3.065 ;
      RECT 1.735 1.635 2.065 2.675 ;
      RECT 0.115 2.145 2.065 2.315 ;
  END
END scs130lp_nor4_lp

MACRO scs130lp_nor4_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.19 0.805 1.86 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 1.19 1.285 1.86 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.58 1.19 1.765 1.86 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.41 0.84 2.725 1.75 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 2.055 2.285 2.845 ;
        RECT 0.09 2.055 2.285 2.225 ;
        RECT 0.09 0.84 2.035 1.01 ;
        RECT 1.825 0.46 2.035 1.01 ;
        RECT 0.635 0.46 0.935 1.01 ;
        RECT 0.09 0.84 0.26 2.225 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.255 -0.085 2.465 0.66 ;
        RECT 1.115 -0.085 1.445 0.6 ;
        RECT 0.245 -0.085 0.455 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 0.475 2.405 0.685 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
END scs130lp_nor4_m

MACRO scs130lp_nor4b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4b_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.095 1.285 1.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.335 1.895 1.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.345 2.355 1.8 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.425 0.595 1.76 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8862 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.865 1.845 3.275 3.075 ;
        RECT 3.065 0.985 3.275 3.075 ;
        RECT 1.455 0.995 3.275 1.165 ;
        RECT 2.355 0.985 3.275 1.165 ;
        RECT 2.355 0.255 2.6 1.165 ;
        RECT 1.455 0.255 1.685 1.165 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.77 -0.085 3.1 0.815 ;
        RECT 1.855 -0.085 2.185 0.825 ;
        RECT 0.79 -0.085 1.24 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 0.9 2.31 1.23 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.36 1.97 2.695 2.14 ;
      RECT 2.525 1.345 2.695 2.14 ;
      RECT 0.36 1.93 0.935 2.14 ;
      RECT 0.765 1.085 0.935 2.14 ;
      RECT 2.525 1.345 2.895 1.675 ;
      RECT 0.36 1.085 0.935 1.255 ;
      RECT 0.36 0.7 0.62 1.255 ;
  END
END scs130lp_nor4b_1

MACRO scs130lp_nor4b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4b_2 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.87 1.21 4.645 1.445 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.4 1.615 5.195 1.785 ;
        RECT 4.815 1.185 5.195 1.785 ;
        RECT 3.4 1.345 3.66 1.785 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.49 1.085 2.88 1.515 ;
        RECT 0.865 1.085 2.88 1.255 ;
        RECT 0.865 1.085 1.065 1.515 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.185 0.355 1.515 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.06 0.87 4.685 1.04 ;
        RECT 4.495 0.265 4.685 1.04 ;
        RECT 1.535 0.745 3.825 0.915 ;
        RECT 3.565 0.255 3.825 1.04 ;
        RECT 3.06 0.745 3.7 1.175 ;
        RECT 1.585 1.805 3.23 1.975 ;
        RECT 3.06 0.745 3.23 1.975 ;
        RECT 1.585 1.805 2.735 2.145 ;
        RECT 2.465 0.255 2.725 0.915 ;
        RECT 1.535 0.255 1.795 0.915 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.855 -0.085 5.185 1.015 ;
        RECT 3.995 -0.085 4.325 0.7 ;
        RECT 2.985 -0.085 3.315 0.575 ;
        RECT 1.965 -0.085 2.295 0.575 ;
        RECT 0.865 -0.085 1.365 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.935 2.455 5.195 3.415 ;
        RECT 3.995 2.455 5.195 2.665 ;
        RECT 0.525 2.72 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.905 2.145 3.235 3.075 ;
      RECT 1.105 2.035 1.41 3.075 ;
      RECT 1.105 2.315 3.235 2.485 ;
      RECT 2.905 2.145 3.815 2.315 ;
      RECT 1.105 2.035 1.415 2.485 ;
      RECT 3.645 2.005 5.185 2.285 ;
      RECT 3.44 2.835 4.755 3.075 ;
      RECT 3.44 2.485 3.77 3.075 ;
      RECT 0.095 1.695 0.355 3.05 ;
      RECT 0.095 1.695 1.415 1.865 ;
      RECT 1.245 1.425 1.415 1.865 ;
      RECT 0.525 0.795 0.695 1.865 ;
      RECT 1.245 1.425 2.32 1.635 ;
      RECT 0.15 0.795 0.695 1.005 ;
      RECT 1.58 2.655 2.735 3.01 ;
  END
END scs130lp_nor4b_2

MACRO scs130lp_nor4b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4b_4 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.96 1.355 9.03 1.525 ;
        RECT 7.735 1.21 9.03 1.525 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.23 1.355 6.625 1.835 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.01 1.315 4.7 1.485 ;
        RECT 3.885 1.21 4.7 1.485 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.325 0.55 1.76 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.6124 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.045 0.255 8.235 1.04 ;
        RECT 7.145 0.87 8.235 1.04 ;
        RECT 4.87 1.005 7.425 1.185 ;
        RECT 7.145 0.255 7.375 1.185 ;
        RECT 6.285 0.255 6.475 1.185 ;
        RECT 5.425 0.255 5.615 1.185 ;
        RECT 3.205 0.84 5.615 1.04 ;
        RECT 1.475 1.665 5.06 1.835 ;
        RECT 4.87 0.84 5.06 1.835 ;
        RECT 4.065 0.255 4.255 1.04 ;
        RECT 1.095 0.965 3.405 1.145 ;
        RECT 3.205 0.255 3.395 1.145 ;
        RECT 2.335 1.665 2.665 2.735 ;
        RECT 1.965 0.255 2.185 1.145 ;
        RECT 1.475 1.665 1.805 2.735 ;
        RECT 1.095 0.255 1.295 1.145 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 8.405 -0.085 8.735 1.04 ;
        RECT 7.545 -0.085 7.875 0.7 ;
        RECT 6.645 -0.085 6.975 0.835 ;
        RECT 5.785 -0.085 6.115 0.835 ;
        RECT 4.425 -0.085 5.255 0.67 ;
        RECT 3.565 -0.085 3.895 0.67 ;
        RECT 2.355 -0.085 3.035 0.785 ;
        RECT 1.465 -0.085 1.795 0.795 ;
        RECT 0.535 -0.085 0.865 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 8.015 2.105 8.345 3.415 ;
        RECT 7.155 2.105 7.485 3.415 ;
        RECT 0.525 2.27 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.515 1.695 8.775 3.075 ;
      RECT 7.655 1.695 7.845 3.075 ;
      RECT 5.005 2.905 6.985 3.075 ;
      RECT 6.795 1.695 6.985 3.075 ;
      RECT 5.9 2.355 6.125 3.075 ;
      RECT 5.005 2.355 5.335 3.075 ;
      RECT 6.795 1.695 8.775 1.925 ;
      RECT 6.295 2.005 6.625 2.735 ;
      RECT 5.505 2.005 5.73 2.735 ;
      RECT 4.115 2.005 4.315 2.735 ;
      RECT 3.195 2.005 3.525 2.735 ;
      RECT 3.195 2.005 6.625 2.185 ;
      RECT 1.095 2.905 4.815 3.075 ;
      RECT 4.485 2.355 4.815 3.075 ;
      RECT 3.695 2.355 3.895 3.075 ;
      RECT 2.835 2.005 3.025 3.075 ;
      RECT 1.975 2.005 2.165 3.075 ;
      RECT 1.095 1.815 1.305 3.075 ;
      RECT 0.095 1.93 0.355 3.075 ;
      RECT 0.095 1.93 0.925 2.1 ;
      RECT 0.72 0.985 0.925 2.1 ;
      RECT 0.72 1.315 2.8 1.485 ;
      RECT 0.105 0.985 0.925 1.155 ;
      RECT 0.105 0.255 0.365 1.155 ;
  END
END scs130lp_nor4b_4

MACRO scs130lp_nor4b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4b_lp 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 0.905 4.675 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.415 1.215 3.745 2.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.215 3.235 2.89 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.485 1.175 0.835 1.845 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6352 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.54 0.265 3.87 0.725 ;
        RECT 1.565 0.865 3.71 1.035 ;
        RECT 3.54 0.265 3.71 1.035 ;
        RECT 1.565 0.44 2.345 3.065 ;
        RECT 1.875 0.265 2.275 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.33 -0.085 4.66 0.725 ;
        RECT 2.665 -0.085 2.995 0.685 ;
        RECT 1.055 -0.085 1.385 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.21 2.025 4.54 3.415 ;
        RECT 0.665 2.025 0.995 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.135 2.025 0.465 3.065 ;
      RECT 0.135 0.265 0.305 3.065 ;
      RECT 1.055 0.825 1.385 1.845 ;
      RECT 0.135 0.825 1.385 0.995 ;
      RECT 0.135 0.265 0.595 0.995 ;
  END
END scs130lp_nor4b_lp

MACRO scs130lp_nor4b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4b_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.84 1.285 2.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.84 2.12 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.38 2.12 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 0.47 0.805 2.12 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4368 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.91 2.5 3.27 2.83 ;
        RECT 3.1 0.84 3.27 2.83 ;
        RECT 1.515 0.84 3.27 1.01 ;
        RECT 2.355 0.45 2.545 1.01 ;
        RECT 1.515 0.45 1.685 1.01 ;
        RECT 1.355 0.45 1.685 0.66 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.725 -0.085 3.055 0.59 ;
        RECT 1.865 -0.085 2.075 0.65 ;
        RECT 0.985 -0.085 1.175 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.015 2.65 1.345 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.625 2.3 0.835 2.79 ;
      RECT 0.185 2.3 2.73 2.47 ;
      RECT 2.56 1.65 2.92 2.32 ;
      RECT 0.185 0.45 0.395 2.47 ;
  END
END scs130lp_nor4b_m

MACRO scs130lp_nor4bb_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4bb_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 1.105 3.215 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.415 1.425 2.745 1.76 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.735 1.425 4.235 1.76 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.205 0.65 2.12 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8421 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.085 2.855 1.255 ;
        RECT 2.555 0.255 2.855 1.255 ;
        RECT 1.525 1.065 1.945 1.255 ;
        RECT 1.71 0.255 1.945 1.255 ;
        RECT 1.21 1.815 1.695 3.075 ;
        RECT 1.525 1.065 1.695 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.08 -0.085 3.75 0.915 ;
        RECT 2.115 -0.085 2.385 0.915 ;
        RECT 1.16 -0.085 1.54 0.895 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.08 2.315 3.41 3.415 ;
        RECT 0.525 2.63 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.875 1.93 3.95 2.145 ;
      RECT 3.385 1.085 3.555 2.145 ;
      RECT 1.875 1.425 2.205 2.145 ;
      RECT 3.385 1.085 4.16 1.255 ;
      RECT 3.92 0.695 4.16 1.255 ;
      RECT 0.095 2.29 0.355 2.92 ;
      RECT 0.095 2.29 1.03 2.46 ;
      RECT 0.82 1.185 1.03 2.46 ;
      RECT 0.82 1.185 1.355 1.515 ;
      RECT 0.82 0.705 0.99 2.46 ;
      RECT 0.43 0.705 0.99 1.035 ;
  END
END scs130lp_nor4bb_1

MACRO scs130lp_nor4bb_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4bb_2 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.195 1.185 6.635 1.515 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.4 1.185 4.715 1.515 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.58 0.885 2.25 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.58 1.42 2.5 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.885 1.065 6.025 1.235 ;
        RECT 5.835 0.255 6.025 1.235 ;
        RECT 4.885 0.84 5.165 1.235 ;
        RECT 4.975 0.255 5.165 1.235 ;
        RECT 3.635 0.84 5.165 1.015 ;
        RECT 2.705 1.675 4.23 1.845 ;
        RECT 3.995 0.84 4.23 1.845 ;
        RECT 2.775 0.995 4.23 1.165 ;
        RECT 3.635 0.255 3.825 1.165 ;
        RECT 2.705 1.675 3.035 2.735 ;
        RECT 2.775 0.255 2.965 1.165 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 6.195 -0.085 6.525 1.015 ;
        RECT 5.335 -0.085 5.665 0.885 ;
        RECT 3.995 -0.085 4.805 0.67 ;
        RECT 3.135 -0.085 3.465 0.825 ;
        RECT 2.275 -0.085 2.605 0.49 ;
        RECT 0.615 -0.085 0.955 1.07 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 5.845 2.025 6.175 3.415 ;
        RECT 0.635 2.67 1.305 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.345 1.685 6.605 3.075 ;
      RECT 5.485 1.685 5.675 3.075 ;
      RECT 4.555 1.685 4.815 2.735 ;
      RECT 4.555 1.685 6.605 1.855 ;
      RECT 3.585 2.905 5.315 3.075 ;
      RECT 4.985 2.025 5.315 3.075 ;
      RECT 3.585 2.355 3.915 3.075 ;
      RECT 2.275 2.905 3.415 3.075 ;
      RECT 3.205 2.015 3.415 3.075 ;
      RECT 2.275 1.755 2.535 3.075 ;
      RECT 4.085 2.015 4.365 2.735 ;
      RECT 3.205 2.015 4.365 2.185 ;
      RECT 0.185 2.605 0.465 2.935 ;
      RECT 0.185 0.865 0.435 2.935 ;
      RECT 2.385 1.335 3.825 1.505 ;
      RECT 0.185 1.24 1.295 1.41 ;
      RECT 1.125 0.66 1.295 1.41 ;
      RECT 2.385 0.66 2.555 1.505 ;
      RECT 1.125 0.66 2.555 0.83 ;
      RECT 1.475 2.67 1.975 3 ;
      RECT 1.805 1 1.975 3 ;
      RECT 1.805 1 2.205 1.6 ;
      RECT 1.475 1 2.205 1.26 ;
  END
END scs130lp_nor4bb_2

MACRO scs130lp_nor4bb_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4bb_4 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.795 1.375 9.495 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.785 1.355 7.475 1.525 ;
        RECT 5.785 1.355 6.205 1.83 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 1.345 1.285 1.76 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.375 0.475 1.76 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.25 1.005 8.965 1.175 ;
        RECT 8.74 0.255 8.965 1.175 ;
        RECT 7.88 0.255 8.07 1.175 ;
        RECT 7.02 0.255 7.21 1.175 ;
        RECT 4.06 0.995 6.35 1.165 ;
        RECT 6.16 0.255 6.35 1.175 ;
        RECT 4.915 0.985 6.35 1.165 ;
        RECT 3.055 1.685 5.615 1.865 ;
        RECT 5.25 0.985 5.615 1.865 ;
        RECT 4.915 0.255 5.105 1.165 ;
        RECT 4.06 0.255 4.245 1.165 ;
        RECT 2.025 0.655 4.245 0.825 ;
        RECT 4.055 0.255 4.245 0.825 ;
        RECT 3.055 0.255 3.385 0.825 ;
        RECT 3.055 1.685 3.285 2.735 ;
        RECT 2.195 1.685 5.615 1.855 ;
        RECT 2.195 1.685 2.385 2.735 ;
        RECT 2.025 0.255 2.365 0.825 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 9.135 -0.085 9.43 1.095 ;
        RECT 8.24 -0.085 8.57 0.835 ;
        RECT 7.38 -0.085 7.71 0.835 ;
        RECT 6.52 -0.085 6.85 0.835 ;
        RECT 5.275 -0.085 5.99 0.815 ;
        RECT 4.415 -0.085 4.745 0.825 ;
        RECT 3.555 -0.085 3.885 0.485 ;
        RECT 2.535 -0.085 2.865 0.485 ;
        RECT 1.525 -0.085 1.855 0.815 ;
        RECT 0.575 -0.085 0.905 0.855 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 8.67 2.27 9 3.415 ;
        RECT 7.81 2.27 8.14 3.415 ;
        RECT 0.575 2.65 0.905 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.17 1.93 9.43 3.075 ;
      RECT 8.31 1.93 8.5 3.075 ;
      RECT 7.445 1.93 7.64 3.075 ;
      RECT 6.585 1.705 6.775 2.715 ;
      RECT 5.655 2.035 5.915 2.715 ;
      RECT 5.655 2.035 6.775 2.205 ;
      RECT 6.515 1.705 6.775 2.205 ;
      RECT 7.445 1.93 9.43 2.1 ;
      RECT 7.445 1.705 7.625 3.075 ;
      RECT 6.515 1.705 7.625 1.875 ;
      RECT 3.845 2.905 7.275 3.075 ;
      RECT 6.945 2.055 7.275 3.075 ;
      RECT 4.705 2.885 7.275 3.075 ;
      RECT 3.845 2.375 4.175 3.075 ;
      RECT 6.085 2.375 6.415 3.075 ;
      RECT 4.705 2.375 5.035 3.075 ;
      RECT 1.695 2.905 3.675 3.075 ;
      RECT 3.455 2.035 3.675 3.075 ;
      RECT 2.555 2.025 2.885 3.075 ;
      RECT 1.695 2.65 2.025 3.075 ;
      RECT 4.345 2.035 4.535 2.735 ;
      RECT 5.205 2.035 5.465 2.715 ;
      RECT 3.455 2.035 5.465 2.205 ;
      RECT 1.005 1.93 1.635 2.14 ;
      RECT 1.455 0.995 1.635 2.14 ;
      RECT 3.72 1.335 5.07 1.515 ;
      RECT 3.72 0.995 3.89 1.515 ;
      RECT 1.075 0.995 1.635 1.175 ;
      RECT 1.075 0.995 3.89 1.165 ;
      RECT 1.075 0.255 1.335 1.175 ;
      RECT 0.145 1.93 0.405 3.075 ;
      RECT 0.145 2.31 2.025 2.48 ;
      RECT 1.82 1.335 2.025 2.48 ;
      RECT 0.145 1.93 0.825 2.48 ;
      RECT 0.645 1.025 0.825 2.48 ;
      RECT 1.82 1.335 3.51 1.515 ;
      RECT 0.145 1.025 0.825 1.195 ;
      RECT 0.145 0.255 0.395 1.195 ;
  END
END scs130lp_nor4bb_4

MACRO scs130lp_nor4bb_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4bb_lp 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 0.825 4.675 1.495 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.165 3.715 1.495 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 1.175 0.835 1.845 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.855 0.825 5.185 1.495 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5202 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.815 3.785 0.985 ;
        RECT 3.455 0.265 3.785 0.985 ;
        RECT 2.105 1.675 2.625 2.005 ;
        RECT 1.565 0.815 2.275 1.78 ;
        RECT 1.565 0.265 2.175 1.78 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.305 -0.085 4.635 0.645 ;
        RECT 2.635 -0.085 2.965 0.635 ;
        RECT 1.055 -0.085 1.385 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.405 2.025 4.735 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.975 1.675 5.595 3.065 ;
      RECT 5.425 0.265 5.595 3.065 ;
      RECT 2.805 1.675 5.595 1.845 ;
      RECT 2.805 1.165 2.975 1.845 ;
      RECT 2.52 1.165 2.975 1.495 ;
      RECT 5.265 0.265 5.595 0.645 ;
      RECT 1.735 2.895 3.715 3.065 ;
      RECT 3.385 2.025 3.715 3.065 ;
      RECT 1.735 2.535 2.065 3.065 ;
      RECT 1.205 2.025 1.535 3.065 ;
      RECT 2.825 2.025 3.155 2.715 ;
      RECT 1.205 2.185 3.155 2.355 ;
      RECT 0.115 2.025 0.365 3.065 ;
      RECT 0.115 0.265 0.285 3.065 ;
      RECT 1.055 0.825 1.385 1.79 ;
      RECT 0.115 0.825 1.385 0.995 ;
      RECT 0.115 0.265 0.595 0.995 ;
  END
END scs130lp_nor4bb_lp

MACRO scs130lp_nor4bb_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_nor4bb_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.48 1.21 2.81 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.01 0.265 2.725 0.64 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 1.155 3.27 2.49 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.505 0.47 2.175 ;
    END
  END DN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.835 2.575 1.025 ;
        RECT 1.31 1.115 2.245 1.285 ;
        RECT 2.075 0.835 2.245 1.285 ;
        RECT 1.095 2.025 1.48 2.235 ;
        RECT 1.31 0.765 1.48 2.235 ;
        RECT 1.115 0.765 1.48 0.975 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.905 -0.085 3.075 0.935 ;
        RECT 1.66 -0.085 1.83 0.935 ;
        RECT 0.725 -0.085 0.935 0.935 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.665 2.115 2.855 3.415 ;
        RECT 0.525 2.705 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.035 2.855 3.64 3.025 ;
      RECT 3.45 0.765 3.64 3.025 ;
      RECT 3.255 0.765 3.64 0.975 ;
      RECT 0.155 2.355 0.345 2.845 ;
      RECT 0.155 2.355 0.82 2.525 ;
      RECT 0.65 1.155 0.82 2.525 ;
      RECT 0.65 1.155 1.13 1.825 ;
      RECT 0.215 1.155 1.13 1.325 ;
      RECT 0.215 0.795 0.545 1.325 ;
  END
END scs130lp_nor4bb_m

MACRO scs130lp_o2111a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111a_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.035 3.755 2.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.715 1.14 3.215 1.825 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 1.14 2.51 1.865 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 0.375 1.855 1.865 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.08 1.36 1.865 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.385 0.67 3.065 ;
        RECT 0.085 0.265 0.355 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.735 -0.085 3.065 0.525 ;
        RECT 0.525 -0.085 0.855 0.57 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.26 2.385 3.59 3.415 ;
        RECT 1.74 2.385 2.34 3.415 ;
        RECT 0.84 2.385 1.135 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.27 0.695 3.53 0.865 ;
      RECT 3.25 0.28 3.53 0.865 ;
      RECT 2.27 0.28 2.565 0.865 ;
      RECT 2.51 2.035 2.8 3.075 ;
      RECT 1.305 2.035 1.57 3.075 ;
      RECT 0.525 2.035 2.8 2.215 ;
      RECT 0.525 0.74 0.795 2.215 ;
      RECT 0.525 0.74 1.375 0.91 ;
      RECT 1.12 0.28 1.375 0.91 ;
  END
END scs130lp_o2111a_0

MACRO scs130lp_o2111a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111a_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.865 1.335 4.235 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.97 1.335 3.695 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 1.345 2.8 1.76 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 0.39 2.305 1.76 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.325 1.415 1.805 1.76 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 0.255 0.365 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.33 -0.085 3.66 0.825 ;
        RECT 0.535 -0.085 0.855 0.905 ;
        RECT 0.535 -0.085 0.805 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.73 1.93 4.09 3.415 ;
        RECT 2.02 2.27 2.76 3.415 ;
        RECT 0.535 2.27 1.49 3.415 ;
        RECT 0.535 1.815 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.56 0.995 4.09 1.165 ;
      RECT 3.83 0.255 4.09 1.165 ;
      RECT 2.56 0.255 3.16 1.165 ;
      RECT 2.93 1.93 3.26 3.075 ;
      RECT 1.66 1.93 1.85 3.075 ;
      RECT 0.975 1.93 3.26 2.1 ;
      RECT 0.975 1.075 1.145 2.1 ;
      RECT 0.535 1.185 1.145 1.515 ;
      RECT 1.23 0.255 1.56 1.245 ;
      RECT 0.975 1.075 1.56 1.245 ;
  END
END scs130lp_o2111a_1

MACRO scs130lp_o2111a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111a_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.885 1.375 4.235 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 1.425 3.715 2.98 ;
        RECT 3.22 1.425 3.715 1.675 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.58 3.01 1.785 ;
        RECT 2.68 1.425 3.01 1.785 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.01 0.36 2.39 1.535 ;
        RECT 2.01 0.36 2.32 1.785 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.475 1.425 1.84 1.785 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.56 0.255 0.805 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.385 -0.085 3.715 0.865 ;
        RECT 0.975 -0.085 1.285 0.885 ;
        RECT 0.095 -0.085 0.39 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.885 1.92 4.215 3.415 ;
        RECT 2.325 2.295 2.655 3.415 ;
        RECT 0.975 2.295 1.735 3.415 ;
        RECT 0.095 1.82 0.39 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.865 1.035 4.215 1.205 ;
      RECT 3.885 0.255 4.215 1.205 ;
      RECT 2.865 0.255 3.195 1.205 ;
      RECT 2.865 1.955 3.195 3.075 ;
      RECT 1.905 1.955 2.155 3.075 ;
      RECT 1.045 1.955 3.195 2.125 ;
      RECT 1.045 1.055 1.305 2.125 ;
      RECT 0.975 1.055 1.305 1.515 ;
      RECT 0.975 1.055 1.575 1.225 ;
      RECT 1.455 0.255 1.805 1.155 ;
      RECT 1.43 1.02 1.805 1.155 ;
  END
END scs130lp_o2111a_2

MACRO scs130lp_o2111a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111a_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.945 1.415 4.78 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.165 1.325 5.495 1.585 ;
        RECT 5.165 1.075 5.335 1.585 ;
        RECT 3.37 1.075 5.335 1.245 ;
        RECT 3.37 1.075 3.775 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.77 1.425 2.375 1.78 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.425 2.985 1.595 ;
        RECT 1.43 1.95 2.735 2.12 ;
        RECT 2.555 1.425 2.735 2.12 ;
        RECT 1.43 1.425 1.6 2.12 ;
        RECT 1.225 1.425 1.6 1.645 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.39 1.605 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.015 1.755 7.595 1.925 ;
        RECT 7.235 1.065 7.595 1.925 ;
        RECT 5.865 1.065 7.595 1.235 ;
        RECT 6.875 1.755 7.065 3.075 ;
        RECT 6.76 0.255 6.95 1.235 ;
        RECT 6.015 1.755 6.205 3.075 ;
        RECT 5.865 0.255 6.09 1.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.12 -0.085 7.45 0.895 ;
        RECT 6.26 -0.085 6.59 0.895 ;
        RECT 5.43 -0.085 5.695 0.93 ;
        RECT 4.5 -0.085 4.83 0.565 ;
        RECT 3.69 -0.085 3.935 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.235 2.095 7.565 3.415 ;
        RECT 6.375 2.095 6.705 3.415 ;
        RECT 5.515 2.105 5.845 3.415 ;
        RECT 4.11 2.62 4.44 3.415 ;
        RECT 2.35 2.64 2.68 3.415 ;
        RECT 1.445 2.63 1.775 3.415 ;
        RECT 0.55 2.155 0.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.01 1.755 5.3 3.075 ;
      RECT 2.85 2.29 3.545 3.075 ;
      RECT 2.905 1.93 3.545 3.075 ;
      RECT 1.945 2.29 2.18 3.075 ;
      RECT 1.05 2.29 1.275 3.075 ;
      RECT 0.12 1.815 0.38 3.075 ;
      RECT 1.945 2.29 3.545 2.47 ;
      RECT 1.05 2.29 3.545 2.46 ;
      RECT 1.05 1.815 1.25 3.075 ;
      RECT 2.905 1.93 5.3 2.1 ;
      RECT 4.97 1.755 5.3 2.1 ;
      RECT 0.12 1.815 1.25 1.985 ;
      RECT 4.97 1.755 5.845 1.925 ;
      RECT 5.675 1.405 5.845 1.925 ;
      RECT 0.56 0.595 0.89 1.985 ;
      RECT 5.675 1.405 7.055 1.585 ;
      RECT 3.35 0.735 5.26 0.905 ;
      RECT 5 0.255 5.26 0.905 ;
      RECT 3.35 0.725 4.33 0.905 ;
      RECT 4.105 0.255 4.33 0.905 ;
      RECT 3.35 0.255 3.52 0.905 ;
      RECT 1.92 0.255 2.25 0.555 ;
      RECT 1.92 0.255 3.52 0.425 ;
      RECT 4.61 2.28 4.84 3.075 ;
      RECT 3.715 2.28 3.94 3.075 ;
      RECT 3.715 2.28 4.84 2.45 ;
      RECT 1.06 1.085 3.18 1.255 ;
      RECT 2.85 0.595 3.18 1.255 ;
      RECT 1.06 0.255 1.25 1.255 ;
      RECT 0.13 0.255 0.39 1.04 ;
      RECT 0.13 0.255 1.25 0.425 ;
      RECT 1.42 0.725 2.68 0.915 ;
      RECT 2.375 0.68 2.68 0.915 ;
      RECT 1.42 0.285 1.75 0.915 ;
  END
END scs130lp_o2111a_4

MACRO scs130lp_o2111a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111a_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.225 0.67 1.895 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.91 1.225 1.315 1.895 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 0.44 1.825 1.895 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.615 2.395 2.15 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.765 3.235 1.085 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.635 2.075 4.205 3.065 ;
        RECT 3.965 0.265 4.205 3.065 ;
        RECT 3.875 0.265 4.205 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.085 -0.085 3.415 0.585 ;
        RECT 0.555 -0.085 0.885 0.695 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.105 2.075 3.435 3.415 ;
        RECT 1.705 2.68 2.035 3.415 ;
        RECT 0.115 2.075 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.575 1.715 2.905 3.065 ;
      RECT 1.175 2.075 1.505 3.065 ;
      RECT 1.175 2.33 2.905 2.5 ;
      RECT 2.575 1.715 3.745 1.885 ;
      RECT 3.415 1.215 3.745 1.885 ;
      RECT 2.575 1.265 2.745 3.065 ;
      RECT 2.175 1.265 2.745 1.435 ;
      RECT 2.175 0.315 2.345 1.435 ;
      RECT 2.175 0.315 2.715 0.585 ;
      RECT 0.125 0.875 1.315 1.045 ;
      RECT 1.065 0.265 1.315 1.045 ;
      RECT 0.125 0.265 0.375 1.045 ;
  END
END scs130lp_o2111a_lp

MACRO scs130lp_o2111a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111a_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.37 1.21 3.685 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 2.92 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.84 2.335 2.215 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.84 1.795 2.12 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.21 1.285 2.12 ;
    END
  END D1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.785 0.67 2.995 ;
        RECT 0.155 0.265 0.365 2.995 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.925 -0.085 3.135 0.545 ;
        RECT 0.585 -0.085 0.795 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.155 2.845 3.485 3.415 ;
        RECT 1.69 2.845 2.02 3.415 ;
        RECT 0.85 2.785 1.06 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.515 0.725 3.565 0.895 ;
      RECT 3.355 0.345 3.565 0.895 ;
      RECT 2.515 0.345 2.705 0.895 ;
      RECT 2.425 2.435 2.635 2.985 ;
      RECT 1.3 2.435 1.51 2.985 ;
      RECT 0.545 2.435 2.635 2.605 ;
      RECT 0.545 0.725 0.715 2.605 ;
      RECT 0.545 0.725 1.32 0.895 ;
      RECT 1.11 0.345 1.32 0.895 ;
  END
END scs130lp_o2111a_m

MACRO scs130lp_o2111ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111ai_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.155 3.275 2.135 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.155 2.765 2.975 ;
        RECT 2.385 1.155 2.765 1.78 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 0.765 1.855 1.78 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 0.375 1.365 1.78 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 0.765 0.865 1.78 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6445 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.095 1.95 2.355 2.985 ;
        RECT 0.155 1.95 2.355 2.12 ;
        RECT 0.575 1.95 0.885 2.985 ;
        RECT 0.155 0.28 0.85 0.595 ;
        RECT 0.155 0.28 0.365 2.12 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.47 -0.085 2.74 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.935 2.315 3.275 3.415 ;
        RECT 1.055 2.305 1.925 3.415 ;
        RECT 0.125 2.305 0.405 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.035 0.78 3.2 0.95 ;
      RECT 2.91 0.28 3.2 0.95 ;
      RECT 2.035 0.28 2.3 0.95 ;
      RECT 1.65 0.28 2.3 0.595 ;
  END
END scs130lp_o2111ai_0

MACRO scs130lp_o2111ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111ai_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.345 3.235 1.755 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.345 2.735 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.345 1.905 1.76 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 0.38 1.365 1.515 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.61 0.84 0.885 1.515 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5288 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.93 2.365 3.075 ;
        RECT 0.95 1.93 2.365 2.1 ;
        RECT 0.95 1.685 1.365 2.1 ;
        RECT 0.95 1.685 1.285 3.075 ;
        RECT 0.11 1.685 1.365 1.925 ;
        RECT 0.11 0.255 0.78 0.67 ;
        RECT 0.11 0.255 0.44 1.925 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.4 -0.085 2.73 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.9 1.925 3.23 3.415 ;
        RECT 1.48 2.27 1.81 3.415 ;
        RECT 0.43 2.095 0.78 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.84 1.005 3.23 1.175 ;
      RECT 2.9 0.255 3.23 1.175 ;
      RECT 1.84 0.255 2.17 1.175 ;
  END
END scs130lp_o2111ai_1

MACRO scs130lp_o2111ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111ai_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.845 1.185 5.675 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.865 1.185 4.675 1.435 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.445 1.185 3.695 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.375 1.99 1.545 ;
        RECT 1.105 1.21 1.775 1.545 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.425 1.75 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.86 1.685 4.19 2.735 ;
        RECT 2.385 1.685 4.19 1.855 ;
        RECT 2.395 1.685 2.575 3.075 ;
        RECT 0.595 1.755 2.575 1.925 ;
        RECT 1.535 1.755 1.725 3.075 ;
        RECT 0.605 0.595 0.935 1.925 ;
        RECT 0.595 1.165 0.865 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.72 -0.085 5.05 0.675 ;
        RECT 3.86 -0.085 4.19 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.72 1.945 5.05 3.415 ;
        RECT 2.755 2.025 3.085 3.415 ;
        RECT 1.895 2.095 2.225 3.415 ;
        RECT 1.035 2.095 1.365 3.415 ;
        RECT 0.175 1.925 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.57 0.845 5.48 1.015 ;
      RECT 5.22 0.255 5.48 1.015 ;
      RECT 4.36 0.255 4.55 1.015 ;
      RECT 2.57 0.775 3.69 1.015 ;
      RECT 3.5 0.255 3.69 1.015 ;
      RECT 5.22 1.605 5.48 3.075 ;
      RECT 3.43 2.905 4.55 3.075 ;
      RECT 4.36 1.605 4.55 3.075 ;
      RECT 3.43 2.025 3.69 3.075 ;
      RECT 4.36 1.605 5.48 1.775 ;
      RECT 1.505 0.255 1.775 0.7 ;
      RECT 3 0.255 3.33 0.605 ;
      RECT 1.505 0.255 3.33 0.425 ;
      RECT 1.945 0.595 2.275 1.205 ;
      RECT 1.115 0.87 2.275 1.04 ;
      RECT 0.175 0.255 0.435 1.04 ;
      RECT 1.115 0.255 1.335 1.04 ;
      RECT 0.175 0.255 1.335 0.425 ;
  END
END scs130lp_o2111ai_2

MACRO scs130lp_o2111ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111ai_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.925 1.375 9.995 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.01 1.355 7.665 1.525 ;
        RECT 7.135 1.205 7.665 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.945 1.355 5.685 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.085 1.325 3.775 1.505 ;
        RECT 3.115 1.155 3.775 1.505 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 1.335 1.875 1.505 ;
        RECT 0.945 1.2 1.685 1.505 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.0362 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.315 1.705 7.645 2.155 ;
        RECT 6.51 1.705 7.645 1.875 ;
        RECT 6.525 1.705 6.715 2.725 ;
        RECT 3.605 1.92 6.715 2.1 ;
        RECT 6.51 1.705 6.715 2.1 ;
        RECT 5.665 1.92 5.855 3.075 ;
        RECT 4.805 1.92 4.995 3.075 ;
        RECT 3.605 1.92 4.13 3.075 ;
        RECT 3.605 1.675 3.775 3.075 ;
        RECT 0.085 1.675 3.775 1.845 ;
        RECT 2.745 1.675 2.935 3.075 ;
        RECT 1.885 1.675 2.075 3.075 ;
        RECT 0.595 0.7 1.685 1.03 ;
        RECT 1.025 1.675 1.215 3.075 ;
        RECT 0.085 0.985 0.775 1.155 ;
        RECT 0.085 0.985 0.355 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.145 -0.085 9.475 0.835 ;
        RECT 8.285 -0.085 8.615 0.835 ;
        RECT 7.065 -0.085 7.395 0.695 ;
        RECT 6.205 -0.085 6.535 0.845 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.555 1.93 9.885 3.415 ;
        RECT 8.695 2.27 9.025 3.415 ;
        RECT 7.835 2.665 8.165 3.415 ;
        RECT 5.165 2.27 5.495 3.415 ;
        RECT 4.3 2.27 4.635 3.415 ;
        RECT 3.105 2.015 3.435 3.415 ;
        RECT 2.245 2.015 2.575 3.415 ;
        RECT 1.385 2.015 1.715 3.415 ;
        RECT 0.525 2.015 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.055 1.015 6.965 1.185 ;
      RECT 7.835 1.005 9.905 1.175 ;
      RECT 9.645 0.255 9.905 1.175 ;
      RECT 7.565 0.255 8.115 1.035 ;
      RECT 6.705 0.865 8.115 1.035 ;
      RECT 5.845 0.255 6.035 1.185 ;
      RECT 4.985 0.595 5.175 1.185 ;
      RECT 4.055 0.655 4.315 1.185 ;
      RECT 8.785 0.255 8.975 1.175 ;
      RECT 6.705 0.255 6.895 1.185 ;
      RECT 9.195 1.93 9.385 3.075 ;
      RECT 8.335 1.93 8.525 3.075 ;
      RECT 6.025 2.895 7.215 3.075 ;
      RECT 6.885 2.325 7.215 3.075 ;
      RECT 6.025 2.27 6.355 3.075 ;
      RECT 6.885 2.325 8.525 2.495 ;
      RECT 8.265 1.93 8.525 2.495 ;
      RECT 6.885 2.045 7.145 3.075 ;
      RECT 8.265 1.93 9.385 2.1 ;
      RECT 5.345 0.255 5.675 0.845 ;
      RECT 4.485 0.255 4.815 0.845 ;
      RECT 2.245 0.255 2.575 0.815 ;
      RECT 2.245 0.255 4.815 0.485 ;
      RECT 2.245 0.255 5.675 0.425 ;
      RECT 1.855 0.985 2.945 1.155 ;
      RECT 2.745 0.655 3.805 0.985 ;
      RECT 1.855 0.255 2.075 1.155 ;
      RECT 0.095 0.255 0.425 0.815 ;
      RECT 0.095 0.255 2.075 0.53 ;
  END
END scs130lp_o2111ai_4

MACRO scs130lp_o2111ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111ai_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.925 1.18 3.255 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.125 1.125 2.745 1.795 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.125 1.905 1.795 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 0.44 1.375 1.585 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.515 0.905 0.835 1.575 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6797 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.86 1.975 2.19 3.065 ;
        RECT 0.78 1.975 2.19 2.145 ;
        RECT 0.78 1.765 1.11 3.065 ;
        RECT 0.125 1.765 1.11 1.935 ;
        RECT 0.125 0.265 0.71 0.725 ;
        RECT 0.125 0.265 0.335 1.935 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.31 -0.085 2.64 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.89 2.025 3.22 3.415 ;
        RECT 1.31 2.325 1.64 3.415 ;
        RECT 0.25 2.115 0.58 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.8 0.775 3.15 0.945 ;
      RECT 2.82 0.265 3.15 0.945 ;
      RECT 1.8 0.265 2.13 0.945 ;
  END
END scs130lp_o2111ai_lp

MACRO scs130lp_o2111ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2111ai_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 2.885 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.315 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.21 1.855 2.12 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 0.47 1.285 2.12 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.495 0.78 0.805 2.12 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4032 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.82 2.32 2.245 2.965 ;
        RECT 0.635 2.32 2.245 2.625 ;
        RECT 0.635 2.32 1.17 2.985 ;
        RECT 0.145 0.27 0.745 0.6 ;
        RECT 0.145 2.32 2.245 2.49 ;
        RECT 0.145 0.27 0.315 2.49 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.25 -0.085 2.46 0.56 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.55 2.845 2.88 3.415 ;
        RECT 1.39 2.805 1.6 3.415 ;
        RECT 0.265 2.785 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.82 0.74 2.89 0.91 ;
      RECT 2.68 0.36 2.89 0.91 ;
      RECT 1.82 0.36 2.03 0.91 ;
  END
END scs130lp_o2111ai_m

MACRO scs130lp_o211a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211a_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 1.12 1.7 1.565 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.96 1.165 2.28 1.835 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.45 1.53 2.765 1.86 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.915 0.775 3.245 1.02 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4985 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.405 1.065 3.075 ;
        RECT 0.085 0.265 0.365 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.745 -0.085 2.005 0.61 ;
        RECT 0.545 -0.085 0.875 0.615 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.505 2.405 2.765 3.415 ;
        RECT 1.245 2.405 1.575 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.935 1.19 3.265 3.075 ;
      RECT 2.065 2.05 2.335 3.075 ;
      RECT 0.545 2.05 3.265 2.235 ;
      RECT 0.545 1.935 1.79 2.235 ;
      RECT 2.575 1.19 3.265 1.36 ;
      RECT 2.575 0.28 2.745 1.36 ;
      RECT 2.575 0.28 3.265 0.605 ;
      RECT 1.255 0.78 2.405 0.95 ;
      RECT 2.175 0.28 2.405 0.95 ;
      RECT 1.255 0.28 1.575 0.95 ;
  END
END scs130lp_o211a_0

MACRO scs130lp_o211a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211a_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.365 1.825 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.365 2.365 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.535 1.365 3.205 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.365 3.755 1.75 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.815 0.86 3.075 ;
        RECT 0.085 0.255 0.415 1 ;
        RECT 0.085 0.255 0.33 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.815 -0.085 2.145 0.515 ;
        RECT 0.585 -0.085 0.915 1.015 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.75 2.26 3.08 3.415 ;
        RECT 1.03 2.26 1.7 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.25 1.92 3.57 3.075 ;
      RECT 2.215 1.92 2.545 3.075 ;
      RECT 1.085 1.92 3.57 2.09 ;
      RECT 1.085 1.025 1.325 2.09 ;
      RECT 0.5 1.185 1.325 1.515 ;
      RECT 3.24 0.255 3.57 1.195 ;
      RECT 1.085 1.025 3.57 1.195 ;
      RECT 1.29 0.685 2.725 0.855 ;
      RECT 2.395 0.255 2.725 0.855 ;
      RECT 1.29 0.255 1.62 0.855 ;
  END
END scs130lp_o211a_1

MACRO scs130lp_o211a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211a_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.025 1.21 2.32 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.815 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.93 1.21 1.285 1.47 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.355 1.575 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.03 1.25 3.485 2.12 ;
        RECT 3.035 1.25 3.225 3.075 ;
        RECT 3.03 1.19 3.22 2.46 ;
        RECT 3.03 0.955 3.2 2.46 ;
        RECT 2.735 0.255 3.065 1.125 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.37 -0.085 3.62 1.055 ;
        RECT 3.235 -0.085 3.62 0.785 ;
        RECT 2.335 -0.085 2.565 1.04 ;
        RECT 1.405 -0.085 1.735 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.395 2.29 3.725 3.415 ;
        RECT 2.195 2.63 2.865 3.415 ;
        RECT 0.715 2.085 1.045 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.215 2.29 1.615 3.075 ;
      RECT 0.265 1.745 0.545 3.075 ;
      RECT 1.215 2.29 2.66 2.46 ;
      RECT 2.49 1.295 2.66 2.46 ;
      RECT 1.215 1.64 1.425 3.075 ;
      RECT 0.525 1.64 1.425 1.915 ;
      RECT 0.525 0.86 0.705 1.915 ;
      RECT 2.49 1.295 2.86 1.625 ;
      RECT 0.095 0.86 0.705 1.04 ;
      RECT 0.095 0.255 0.425 1.04 ;
      RECT 0.885 0.87 2.165 1.04 ;
      RECT 1.905 0.27 2.165 1.04 ;
      RECT 0.885 0.27 1.215 1.04 ;
  END
END scs130lp_o211a_2

MACRO scs130lp_o211a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211a_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.315 1.085 6.635 1.76 ;
        RECT 4.83 1.085 6.635 1.255 ;
        RECT 4.67 1.195 5 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.21 1.425 6.145 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.93 4.46 2.1 ;
        RECT 4.13 1.345 4.46 2.1 ;
        RECT 2.545 1.405 3.275 2.1 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.445 1.405 3.92 1.76 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.845 1.755 2.035 3.075 ;
        RECT 0.085 1.755 2.035 1.925 ;
        RECT 0.085 1.045 1.655 1.215 ;
        RECT 1.455 0.255 1.655 1.215 ;
        RECT 0.985 1.755 1.165 3.075 ;
        RECT 0.595 0.255 0.785 1.215 ;
        RECT 0.085 1.045 0.37 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.835 -0.085 6.025 0.575 ;
        RECT 4.835 -0.085 5.165 0.575 ;
        RECT 1.85 -0.085 2.085 0.94 ;
        RECT 0.955 -0.085 1.285 0.875 ;
        RECT 0.095 -0.085 0.425 0.875 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 6.195 1.93 6.525 3.415 ;
        RECT 4.47 2.61 4.735 3.415 ;
        RECT 3.465 2.61 3.795 3.415 ;
        RECT 2.205 2.61 2.535 3.415 ;
        RECT 1.345 2.095 1.675 3.415 ;
        RECT 0.485 2.095 0.815 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.365 0.635 4.66 1.025 ;
      RECT 4.365 0.745 6.525 0.915 ;
      RECT 6.195 0.255 6.525 0.915 ;
      RECT 2.335 0.255 2.665 0.895 ;
      RECT 2.335 0.635 4.665 0.805 ;
      RECT 5.335 0.255 5.665 0.915 ;
      RECT 4.395 0.255 4.665 0.915 ;
      RECT 4.905 2.78 6.025 3.075 ;
      RECT 5.835 1.93 6.025 3.075 ;
      RECT 3.965 2.27 4.3 3.075 ;
      RECT 2.705 2.27 3.295 3.075 ;
      RECT 5.335 1.93 5.665 2.61 ;
      RECT 2.205 2.27 5.665 2.44 ;
      RECT 2.205 1.065 2.375 2.44 ;
      RECT 0.54 1.385 2.375 1.585 ;
      RECT 2.205 1.065 3.7 1.235 ;
      RECT 3.37 0.975 3.7 1.235 ;
      RECT 2.845 0.255 4.225 0.465 ;
  END
END scs130lp_o211a_4

MACRO scs130lp_o211a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211a_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 1.44 0.57 2.14 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.78 1.44 1.42 2.14 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.59 1.55 1.87 2.14 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.345 3.235 1.78 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.475 0.265 3.725 3.065 ;
        RECT 3.395 0.265 3.725 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.575 -0.085 2.905 0.615 ;
        RECT 0.625 -0.085 0.955 0.93 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.865 2.025 3.195 3.415 ;
        RECT 1.665 2.66 1.995 3.415 ;
        RECT 0.115 2.31 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.175 2.075 2.635 3.065 ;
      RECT 1.135 2.31 1.465 3.065 ;
      RECT 1.135 2.31 2.635 2.48 ;
      RECT 2.175 0.795 2.345 3.065 ;
      RECT 1.955 0.7 2.285 1.16 ;
      RECT 1.955 0.795 3.21 1.125 ;
      RECT 0.115 1.1 1.41 1.27 ;
      RECT 1.135 0.7 1.465 1.16 ;
      RECT 0.115 0.85 0.365 1.27 ;
  END
END scs130lp_o211a_lp

MACRO scs130lp_o211a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211a_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 0.985 1.415 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.985 2.04 1.495 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 2.515 2.4 3.025 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.805 0.84 3.205 1.51 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 2.025 0.75 2.86 ;
        RECT 0.095 0.47 0.425 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.475 -0.085 1.805 0.455 ;
        RECT 0.605 -0.085 0.795 0.74 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.58 2.045 2.75 3.415 ;
        RECT 2.42 2.045 2.75 2.255 ;
        RECT 0.945 2.025 1.275 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.93 1.695 3.12 2.165 ;
      RECT 1.895 1.675 2.105 2.165 ;
      RECT 1.895 1.695 3.12 1.865 ;
      RECT 0.625 1.675 2.625 1.845 ;
      RECT 2.455 0.33 2.625 1.865 ;
      RECT 0.625 1.025 0.795 1.845 ;
      RECT 2.455 0.33 3.045 0.66 ;
      RECT 1.105 0.635 2.255 0.805 ;
      RECT 2.045 0.355 2.255 0.805 ;
      RECT 1.105 0.355 1.295 0.805 ;
  END
END scs130lp_o211a_m

MACRO scs130lp_o211ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211ai_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.08 0.575 1.85 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 1.08 1.295 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.08 1.84 1.78 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.4 0.785 2.795 1.78 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4601 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.22 1.95 2.795 2.985 ;
        RECT 2.01 0.28 2.46 0.615 ;
        RECT 2.01 0.28 2.22 2.135 ;
        RECT 0.99 1.95 2.795 2.135 ;
        RECT 0.99 1.95 1.29 2.985 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.57 -0.085 1.24 0.57 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.46 2.305 2.05 3.415 ;
        RECT 0.2 2.305 0.53 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.14 0.74 1.67 0.91 ;
      RECT 1.41 0.28 1.67 0.91 ;
      RECT 0.14 0.28 0.4 0.91 ;
  END
END scs130lp_o211ai_0

MACRO scs130lp_o211ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211ai_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.185 0.435 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.185 1.09 1.515 ;
        RECT 0.605 1.185 0.845 2.86 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.3 1.345 1.795 1.78 ;
        RECT 1.57 0.39 1.795 1.78 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.965 1.295 2.3 1.78 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.7619 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 1.95 2.78 3.075 ;
        RECT 2.47 0.255 2.78 3.075 ;
        RECT 1.965 0.255 2.78 1.095 ;
        RECT 1.015 1.95 2.78 2.12 ;
        RECT 1.015 1.95 1.28 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.595 -0.085 0.925 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.48 2.29 1.81 3.415 ;
        RECT 0.095 1.92 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.095 0.845 1.4 1.015 ;
      RECT 1.125 0.255 1.4 1.015 ;
      RECT 0.095 0.255 0.425 1.015 ;
  END
END scs130lp_o211ai_1

MACRO scs130lp_o211ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211ai_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.56 1.42 4.715 1.59 ;
        RECT 4.115 1.21 4.715 1.59 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.42 3.28 1.59 ;
        RECT 2.075 1.195 2.735 1.59 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.21 1.905 1.525 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.285 0.445 1.75 ;
        RECT 0.085 1.21 0.385 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.825 1.76 3.155 2.735 ;
        RECT 0.615 1.76 3.155 1.93 ;
        RECT 1.475 1.76 1.665 3.075 ;
        RECT 0.615 0.595 0.875 1.93 ;
        RECT 0.615 0.595 0.805 3.075 ;
        RECT 0.545 0.595 0.875 1.145 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.115 -0.085 4.445 1.04 ;
        RECT 3.255 -0.085 3.585 0.91 ;
        RECT 2.395 -0.085 2.725 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.685 2.1 4.015 3.415 ;
        RECT 1.835 2.1 2.165 3.415 ;
        RECT 0.975 2.1 1.305 3.415 ;
        RECT 0.115 1.92 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.185 1.76 4.445 3.075 ;
      RECT 2.395 2.905 3.515 3.075 ;
      RECT 3.325 1.76 3.515 3.075 ;
      RECT 2.395 2.1 2.655 3.075 ;
      RECT 3.325 1.76 4.445 1.93 ;
      RECT 2.905 1.08 3.945 1.25 ;
      RECT 3.755 0.255 3.945 1.25 ;
      RECT 2.905 0.255 3.085 1.25 ;
      RECT 1.405 0.815 3.085 1.025 ;
      RECT 2.895 0.255 3.085 1.025 ;
      RECT 1.045 0.255 1.235 1.04 ;
      RECT 0.095 0.255 0.375 1.04 ;
      RECT 1.045 0.255 2.165 0.645 ;
      RECT 0.095 0.255 2.165 0.425 ;
  END
END scs130lp_o211ai_2

MACRO scs130lp_o211ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211ai_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.925 3.78 2.12 ;
        RECT 3.5 1.345 3.78 2.12 ;
        RECT 1.115 1.345 1.56 2.12 ;
        RECT 0.21 1.345 1.56 1.63 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.855 1.425 3.33 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.955 1.93 7.72 2.1 ;
        RECT 7.39 1.425 7.72 2.1 ;
        RECT 4.955 1.345 5.125 2.1 ;
        RECT 3.95 1.345 5.125 1.76 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.355 1.425 7.045 1.76 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.5872 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.9 2.27 8.07 2.505 ;
        RECT 7.89 1.075 8.07 2.505 ;
        RECT 5.675 1.075 8.07 1.255 ;
        RECT 7.145 2.27 7.335 3.075 ;
        RECT 5.675 0.965 7.025 1.255 ;
        RECT 5.9 2.27 6.135 3.075 ;
        RECT 4.215 2.27 8.07 2.44 ;
        RECT 5.085 2.27 5.31 3.075 ;
        RECT 4.215 1.93 4.425 2.44 ;
        RECT 4.205 2.29 4.415 3.075 ;
        RECT 2.025 2.29 4.415 2.51 ;
        RECT 2.025 2.29 2.235 2.63 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 3.255 -0.085 3.585 0.825 ;
        RECT 2.395 -0.085 2.725 0.825 ;
        RECT 1.535 -0.085 1.865 0.805 ;
        RECT 0.675 -0.085 1.005 0.825 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.505 2.675 7.835 3.415 ;
        RECT 6.305 2.675 6.975 3.415 ;
        RECT 5.48 2.61 5.73 3.415 ;
        RECT 4.585 2.61 4.915 3.415 ;
        RECT 3.705 2.68 4.035 3.415 ;
        RECT 1.105 2.69 1.435 3.415 ;
        RECT 0.245 1.815 0.535 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.305 0.995 4.915 1.175 ;
      RECT 4.655 0.625 4.915 1.175 ;
      RECT 3.755 0.255 3.985 1.175 ;
      RECT 2.895 0.255 3.085 1.175 ;
      RECT 2.035 0.255 2.225 1.175 ;
      RECT 1.175 0.255 1.365 1.175 ;
      RECT 0.305 0.255 0.505 1.175 ;
      RECT 7.715 0.365 8.045 0.905 ;
      RECT 4.655 0.625 8.045 0.795 ;
      RECT 4.155 0.265 4.485 0.825 ;
      RECT 4.155 0.265 7.535 0.455 ;
      RECT 1.605 2.81 3.525 3.075 ;
      RECT 3.315 2.68 3.525 3.075 ;
      RECT 0.705 1.815 0.925 3.075 ;
      RECT 1.605 2.29 1.805 3.075 ;
      RECT 0.705 2.29 1.805 2.52 ;
  END
END scs130lp_o211ai_4

MACRO scs130lp_o211ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211ai_lp 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.17 0.625 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.925 1.17 1.315 1.84 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.17 1.825 1.84 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.11 2.395 1.78 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7247 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.29 2.02 2.755 3.065 ;
        RECT 2.585 0.265 2.755 3.065 ;
        RECT 2.01 0.265 2.755 0.725 ;
        RECT 1.19 2.02 2.755 2.19 ;
        RECT 1.19 2.02 1.52 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.68 -0.085 1.01 0.64 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.72 2.37 2.05 3.415 ;
        RECT 0.13 2.025 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.17 0.82 1.52 0.99 ;
      RECT 1.19 0.265 1.52 0.99 ;
      RECT 0.17 0.265 0.5 0.99 ;
  END
END scs130lp_o211ai_lp

MACRO scs130lp_o211ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o211ai_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.47 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.77 1.015 1.285 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.31 1.705 1.765 2.215 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.85 0.84 2.245 1.015 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3402 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.58 2.245 2.985 ;
        RECT 1.945 1.195 2.115 2.665 ;
        RECT 1.5 0.33 2.065 0.66 ;
        RECT 1.135 2.495 2.245 2.665 ;
        RECT 1.5 1.195 2.115 1.365 ;
        RECT 1.5 0.33 1.67 1.365 ;
        RECT 1.135 2.495 1.345 2.985 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.555 -0.085 0.885 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.525 2.845 1.855 3.415 ;
        RECT 0.285 2.845 0.615 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.165 0.665 1.275 0.835 ;
      RECT 1.065 0.345 1.275 0.835 ;
      RECT 0.165 0.345 0.375 0.835 ;
  END
END scs130lp_o211ai_m

MACRO scs130lp_o21a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21a_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.01 1.175 2.555 2.225 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.175 1.84 2.97 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 1.125 1.365 1.795 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.395 0.565 3.075 ;
        RECT 0.085 0.275 0.4 0.605 ;
        RECT 0.085 0.275 0.335 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.935 -0.085 2.205 0.665 ;
        RECT 0.57 -0.085 0.855 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.02 2.395 2.35 3.415 ;
        RECT 0.735 2.395 1.005 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.515 0.835 2.665 1.005 ;
      RECT 2.375 0.335 2.665 1.005 ;
      RECT 1.515 0.335 1.765 1.005 ;
      RECT 1.175 2.045 1.425 3.075 ;
      RECT 0.505 2.045 1.425 2.215 ;
      RECT 0.505 0.775 0.755 2.215 ;
      RECT 0.505 0.775 1.345 0.955 ;
      RECT 1.105 0.335 1.345 0.955 ;
  END
END scs130lp_o21a_0

MACRO scs130lp_o21a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21a_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.375 2.795 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.425 2.255 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.075 1.425 1.415 1.76 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.695 0.545 3.075 ;
        RECT 0.085 0.255 0.355 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.955 -0.085 2.285 0.855 ;
        RECT 0.525 -0.085 0.855 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.435 1.93 2.765 3.415 ;
        RECT 0.715 2.27 1.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.515 1.025 2.765 1.195 ;
      RECT 2.455 0.255 2.765 1.195 ;
      RECT 1.515 0.255 1.785 1.195 ;
      RECT 1.605 1.93 1.935 3.075 ;
      RECT 0.735 1.93 1.935 2.1 ;
      RECT 0.735 1.085 0.905 2.1 ;
      RECT 0.525 1.085 0.905 1.515 ;
      RECT 0.525 1.085 1.345 1.255 ;
      RECT 1.045 0.255 1.345 1.255 ;
  END
END scs130lp_o21a_1

MACRO scs130lp_o21a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21a_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.375 3.275 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.375 2.735 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.485 1.415 1.895 1.75 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.565 0.255 0.815 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.385 -0.085 2.715 0.865 ;
        RECT 0.985 -0.085 1.315 0.905 ;
        RECT 0.125 -0.085 0.395 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.835 1.92 3.165 3.415 ;
        RECT 0.985 2.26 1.835 3.415 ;
        RECT 0.125 1.815 0.395 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.97 1.035 3.165 1.205 ;
      RECT 2.885 0.255 3.165 1.205 ;
      RECT 1.97 0.255 2.215 1.205 ;
      RECT 2.005 1.92 2.265 3.075 ;
      RECT 1.145 1.92 2.265 2.09 ;
      RECT 1.145 1.075 1.315 2.09 ;
      RECT 0.985 1.075 1.315 1.52 ;
      RECT 0.985 1.075 1.8 1.245 ;
      RECT 1.505 0.255 1.8 1.245 ;
  END
END scs130lp_o21a_2

MACRO scs130lp_o21a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21a_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.955 1.425 5.43 1.645 ;
        RECT 3.745 2.31 5.125 2.5 ;
        RECT 4.955 1.425 5.125 2.5 ;
        RECT 3.745 1.425 3.915 2.5 ;
        RECT 3.585 1.425 3.915 1.675 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 1.425 4.775 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 1.425 3.185 1.76 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.825 1.755 2.005 3.075 ;
        RECT 0.085 1.755 2.005 1.925 ;
        RECT 0.085 1.055 1.695 1.225 ;
        RECT 1.505 0.255 1.695 1.225 ;
        RECT 0.965 1.755 1.155 3.075 ;
        RECT 0.645 0.255 0.835 1.225 ;
        RECT 0.085 1.055 0.35 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.795 -0.085 5.125 0.915 ;
        RECT 3.925 -0.085 4.265 0.565 ;
        RECT 1.865 -0.085 2.195 0.905 ;
        RECT 1.005 -0.085 1.335 0.885 ;
        RECT 0.145 -0.085 0.475 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.295 1.815 5.555 3.415 ;
        RECT 3.045 2.805 3.815 3.415 ;
        RECT 3.245 1.925 3.575 3.415 ;
        RECT 2.185 2.27 2.515 3.415 ;
        RECT 1.325 2.095 1.655 3.415 ;
        RECT 0.465 2.095 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.435 1.085 5.555 1.255 ;
      RECT 5.295 0.305 5.555 1.255 ;
      RECT 4.435 0.305 4.625 1.255 ;
      RECT 3.425 0.735 4.625 0.905 ;
      RECT 2.415 0.255 2.745 0.895 ;
      RECT 3.425 0.255 3.755 0.905 ;
      RECT 2.415 0.255 3.755 0.425 ;
      RECT 2.685 1.93 2.875 3.075 ;
      RECT 4.085 1.93 4.695 2.14 ;
      RECT 2.175 1.93 2.875 2.1 ;
      RECT 4.085 1.075 4.265 2.14 ;
      RECT 2.175 1.075 2.345 2.1 ;
      RECT 0.52 1.395 2.345 1.585 ;
      RECT 2.175 1.075 4.265 1.245 ;
      RECT 2.915 0.595 3.245 1.245 ;
      RECT 3.995 2.67 5.065 3 ;
  END
END scs130lp_o21a_4

MACRO scs130lp_o21a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21a_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.175 0.55 1.845 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.87 1.18 1.315 2.89 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.175 1.825 1.505 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 2.105 3.245 2.275 ;
        RECT 2.915 0.295 3.245 2.275 ;
        RECT 2.555 2.105 2.885 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.125 -0.085 2.455 0.645 ;
        RECT 0.625 -0.085 0.875 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.025 2.035 2.355 3.415 ;
        RECT 0.175 2.025 0.505 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.495 1.685 1.825 3.065 ;
      RECT 1.495 1.685 2.175 1.855 ;
      RECT 2.005 0.825 2.175 1.855 ;
      RECT 2.355 0.825 2.685 1.495 ;
      RECT 1.565 0.825 2.685 0.995 ;
      RECT 1.565 0.265 1.895 0.995 ;
      RECT 0.115 0.825 1.385 0.995 ;
      RECT 1.055 0.265 1.385 0.995 ;
      RECT 0.115 0.265 0.445 0.995 ;
  END
END scs130lp_o21a_lp

MACRO scs130lp_o21a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21a_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.42 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.8 2.49 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 1.21 1.285 2.12 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.715 0.715 2.925 ;
        RECT 0.155 0.265 0.365 0.595 ;
        RECT 0.155 0.265 0.325 2.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.965 -0.085 2.175 0.68 ;
        RECT 0.585 -0.085 0.795 0.555 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.035 2.845 2.365 3.415 ;
        RECT 0.895 2.785 1.065 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.535 0.86 2.605 1.03 ;
      RECT 2.395 0.48 2.605 1.03 ;
      RECT 1.535 0.48 1.745 1.03 ;
      RECT 1.245 2.715 1.575 2.925 ;
      RECT 1.245 2.3 1.415 2.925 ;
      RECT 0.505 2.3 1.415 2.47 ;
      RECT 0.505 0.775 0.675 2.47 ;
      RECT 0.505 0.775 1.315 0.945 ;
      RECT 1.105 0.48 1.315 0.945 ;
  END
END scs130lp_o21a_m

MACRO scs130lp_o21ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ai_0 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.015 0.455 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.1 0.92 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.45 1.47 1.835 2.15 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2905 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.1 1.12 1.775 1.29 ;
        RECT 1.49 0.28 1.775 1.29 ;
        RECT 1.015 2.32 1.335 3.075 ;
        RECT 1.1 2.28 1.335 3.075 ;
        RECT 1.1 1.12 1.27 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.585 -0.085 0.915 0.505 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.505 2.395 1.775 3.415 ;
        RECT 0.195 2.395 0.525 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.155 0.675 1.32 0.845 ;
      RECT 1.085 0.28 1.32 0.845 ;
      RECT 0.155 0.28 0.415 0.845 ;
  END
END scs130lp_o21ai_0

MACRO scs130lp_o21ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ai_1 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.415 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.585 1.345 1.02 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.315 1.835 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7896 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.19 0.975 1.825 1.145 ;
        RECT 1.565 0.255 1.825 1.145 ;
        RECT 0.94 1.92 1.36 3.075 ;
        RECT 1.19 0.975 1.36 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.565 -0.085 0.895 0.465 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.53 1.92 1.825 3.415 ;
        RECT 0.105 1.92 0.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.105 0.635 1.02 1.04 ;
      RECT 0.105 0.635 1.395 0.805 ;
      RECT 1.065 0.255 1.395 0.805 ;
      RECT 0.105 0.265 0.375 1.04 ;
  END
END scs130lp_o21ai_1

MACRO scs130lp_o21ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ai_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.245 1.345 2.355 1.75 ;
        RECT 0.125 1.695 1.415 1.865 ;
        RECT 0.125 1.375 0.455 1.865 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.185 1.025 1.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.21 3.265 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9408 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.5 1.92 2.735 3.075 ;
        RECT 2.525 0.595 2.735 3.075 ;
        RECT 1 2.035 2.735 2.205 ;
        RECT 1.595 1.92 2.735 2.205 ;
        RECT 1 2.035 1.3 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.535 -0.085 1.865 0.825 ;
        RECT 0.54 -0.085 0.87 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.905 1.92 3.215 3.415 ;
        RECT 2 2.375 2.33 3.415 ;
        RECT 0.11 2.035 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.195 1.005 2.355 1.175 ;
      RECT 2.035 0.255 2.355 1.175 ;
      RECT 2.905 0.255 3.215 1.04 ;
      RECT 1.04 0.255 1.365 1.015 ;
      RECT 0.11 0.845 1.365 1.015 ;
      RECT 0.11 0.255 0.37 1.015 ;
      RECT 2.035 0.255 3.215 0.425 ;
      RECT 0.61 2.905 1.805 3.075 ;
      RECT 1.475 2.375 1.805 3.075 ;
      RECT 0.61 2.035 0.83 3.075 ;
  END
END scs130lp_o21ai_2

MACRO scs130lp_o21ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ai_4 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.445 1.075 3.695 1.515 ;
        RECT 1.42 1.075 3.695 1.245 ;
        RECT 0.125 1.21 1.825 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 1.425 3.275 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.905 1.21 5.255 1.435 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8816 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.425 0.7 5.67 1.925 ;
        RECT 3.865 1.605 5.67 1.925 ;
        RECT 4.1 0.7 5.67 1.03 ;
        RECT 4.96 1.605 5.15 3.075 ;
        RECT 4.08 1.605 4.29 3.075 ;
        RECT 1.84 1.93 4.29 2.1 ;
        RECT 3.445 1.755 4.29 2.1 ;
        RECT 2.7 1.93 3.03 2.735 ;
        RECT 1.84 1.93 2.17 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 3.13 -0.085 3.46 0.565 ;
        RECT 2.27 -0.085 2.6 0.565 ;
        RECT 1.41 -0.085 1.74 0.565 ;
        RECT 0.55 -0.085 0.88 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.32 2.105 5.65 3.415 ;
        RECT 4.46 2.095 4.79 3.415 ;
        RECT 3.58 2.27 3.91 3.415 ;
        RECT 0.98 2.095 1.31 3.415 ;
        RECT 0.12 1.815 0.405 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.12 0.87 1.25 1.04 ;
      RECT 3.63 0.255 3.93 0.905 ;
      RECT 1.05 0.735 3.93 0.905 ;
      RECT 0.12 0.255 0.38 1.04 ;
      RECT 2.77 0.255 2.96 0.905 ;
      RECT 1.91 0.255 2.1 0.905 ;
      RECT 1.05 0.255 1.24 1.04 ;
      RECT 3.63 0.255 5.65 0.53 ;
      RECT 1.48 2.905 3.41 3.075 ;
      RECT 3.2 2.27 3.41 3.075 ;
      RECT 0.575 1.755 0.81 3.075 ;
      RECT 2.34 2.27 2.53 3.075 ;
      RECT 1.48 1.755 1.67 3.075 ;
      RECT 0.575 1.755 1.67 1.925 ;
  END
END scs130lp_o21ai_4

MACRO scs130lp_o21ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ai_lp 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.125 0.835 1.795 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.125 1.345 1.795 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.125 1.915 1.795 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4733 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.24 1.975 2.265 2.145 ;
        RECT 2.095 0.265 2.265 2.145 ;
        RECT 1.83 0.265 2.265 0.725 ;
        RECT 1.24 1.975 1.57 3.065 ;
        RECT 1.085 2.29 1.57 2.89 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 0.81 -0.085 1.14 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.81 2.325 2.14 3.415 ;
        RECT 0.22 2.025 0.55 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.3 0.775 1.65 0.945 ;
      RECT 1.32 0.265 1.65 0.945 ;
      RECT 0.3 0.265 0.63 0.945 ;
  END
END scs130lp_o21ai_lp

MACRO scs130lp_o21ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ai_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.035 0.455 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 2.69 1.285 3 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.08 1.47 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2835 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.93 1.82 2.1 ;
        RECT 1.65 0.425 1.82 2.1 ;
        RECT 1.405 0.425 1.82 0.635 ;
        RECT 0.635 1.93 1.285 2.48 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 0.525 -0.085 0.855 0.505 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.485 2.28 1.695 3.415 ;
        RECT 0.095 2.34 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.155 0.685 1.225 0.855 ;
      RECT 1.035 0.365 1.225 0.855 ;
      RECT 0.155 0.365 0.345 0.855 ;
  END
END scs130lp_o21ai_m

MACRO scs130lp_o21ba_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ba_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.015 1.13 3.54 2.215 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.13 2.845 2.205 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.995 0.765 1.305 1.435 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.28 0.465 0.61 ;
        RECT 0.085 1.975 0.355 2.935 ;
        RECT 0.085 0.28 0.335 2.935 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.935 -0.085 3.2 0.61 ;
        RECT 0.635 -0.085 1.305 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.15 2.415 3.48 3.415 ;
        RECT 1.88 2.805 2.21 3.415 ;
        RECT 0.525 1.965 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.505 0.78 3.66 0.96 ;
      RECT 3.37 0.28 3.66 0.96 ;
      RECT 2.505 0.28 2.765 0.96 ;
      RECT 2.38 2.395 2.66 3.075 ;
      RECT 0.975 2.465 2.66 2.635 ;
      RECT 2.1 2.395 2.66 2.635 ;
      RECT 0.975 1.625 1.145 2.635 ;
      RECT 2.1 0.28 2.335 2.635 ;
      RECT 0.505 1.625 1.145 1.795 ;
      RECT 0.505 1.125 0.755 1.795 ;
      RECT 1.315 1.965 1.75 2.295 ;
      RECT 1.475 0.865 1.75 2.295 ;
      RECT 1.475 0.865 1.93 1.535 ;
      RECT 1.475 0.28 1.735 2.295 ;
  END
END scs130lp_o21ba_0

MACRO scs130lp_o21ba_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ba_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.375 3.755 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.48 1.425 3.215 1.75 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.21 1.305 1.75 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5733 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.815 0.575 3.075 ;
        RECT 0.085 0.255 0.385 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.905 -0.085 3.235 0.865 ;
        RECT 0.555 -0.085 0.915 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.405 1.92 3.735 3.415 ;
        RECT 2.015 2.27 2.345 3.415 ;
        RECT 0.745 1.925 1.255 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.48 1.035 3.735 1.205 ;
      RECT 3.405 0.255 3.735 1.205 ;
      RECT 2.48 0.255 2.715 1.205 ;
      RECT 2.525 1.925 2.795 3.075 ;
      RECT 2.075 1.925 2.795 2.1 ;
      RECT 2.075 0.255 2.31 2.1 ;
      RECT 0.565 1.22 0.935 1.55 ;
      RECT 0.765 0.87 0.935 1.55 ;
      RECT 0.765 0.87 1.305 1.04 ;
      RECT 1.135 0.255 1.305 1.04 ;
      RECT 1.135 0.255 2.31 0.425 ;
      RECT 1.425 1.925 1.755 2.21 ;
      RECT 1.475 0.86 1.755 2.21 ;
      RECT 1.475 0.86 1.905 1.55 ;
  END
END scs130lp_o21ba_1

MACRO scs130lp_o21ba_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ba_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.21 3.755 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.785 1.21 3.215 2.605 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.21 0.895 1.75 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 1.85 1.67 2.12 ;
        RECT 1.065 0.255 1.315 2.12 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.935 -0.085 3.265 0.485 ;
        RECT 1.485 -0.085 1.815 0.835 ;
        RECT 0.53 -0.085 0.895 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.385 1.92 3.7 3.415 ;
        RECT 1.84 2.63 2.17 3.415 ;
        RECT 0.91 2.63 1.24 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.375 0.655 3.705 1.04 ;
      RECT 3.435 0.255 3.705 1.04 ;
      RECT 2.435 0.655 3.705 0.835 ;
      RECT 2.435 0.255 2.765 0.835 ;
      RECT 2.405 1.855 2.615 3.075 ;
      RECT 2.435 1.005 2.615 3.075 ;
      RECT 1.485 1.005 1.795 1.515 ;
      RECT 1.485 1.005 2.615 1.175 ;
      RECT 2.005 0.255 2.265 1.175 ;
      RECT 0.085 2.29 2.235 2.46 ;
      RECT 2.005 1.345 2.235 2.46 ;
      RECT 0.085 1.92 0.595 2.46 ;
      RECT 0.085 0.7 0.27 2.46 ;
      RECT 2.005 1.345 2.265 1.675 ;
      RECT 0.085 0.7 0.36 1.03 ;
  END
END scs130lp_o21ba_2

MACRO scs130lp_o21ba_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ba_4 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.435 1.415 5.86 1.645 ;
        RECT 4.075 2.31 5.605 2.5 ;
        RECT 5.435 1.415 5.605 2.5 ;
        RECT 4.075 1.415 4.345 2.5 ;
        RECT 4.015 1.415 4.345 1.675 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.92 1.415 5.25 1.76 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.43 1.2 0.865 1.75 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.93 2.255 2.26 ;
        RECT 1.035 1.075 2.145 1.245 ;
        RECT 1.955 0.255 2.145 1.245 ;
        RECT 1.035 0.255 1.285 1.245 ;
        RECT 0.625 1.92 1.205 2.26 ;
        RECT 1.035 0.255 1.205 2.26 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.225 -0.085 5.555 0.905 ;
        RECT 4.355 -0.085 4.695 0.555 ;
        RECT 2.315 -0.085 2.645 0.905 ;
        RECT 1.455 -0.085 1.785 0.905 ;
        RECT 0.595 -0.085 0.865 1.03 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.775 1.815 6.025 3.415 ;
        RECT 3.595 2.785 4.265 3.415 ;
        RECT 3.595 1.815 3.905 3.415 ;
        RECT 2.36 2.78 3.035 3.415 ;
        RECT 2.765 2.115 3.035 3.415 ;
        RECT 1.495 2.78 1.825 3.415 ;
        RECT 0.635 2.78 0.965 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.865 1.075 6.005 1.245 ;
      RECT 5.735 0.305 6.005 1.245 ;
      RECT 4.865 0.295 5.055 1.245 ;
      RECT 2.835 0.265 3.175 0.905 ;
      RECT 3.855 0.725 5.055 0.895 ;
      RECT 3.855 0.265 4.185 0.895 ;
      RECT 2.835 0.265 4.185 0.435 ;
      RECT 3.205 1.075 3.425 3.075 ;
      RECT 4.525 1.93 5.125 2.14 ;
      RECT 4.525 1.075 4.695 2.14 ;
      RECT 1.375 1.415 2.485 1.605 ;
      RECT 2.315 1.075 2.485 1.605 ;
      RECT 2.315 1.075 4.695 1.245 ;
      RECT 3.345 0.605 3.675 1.245 ;
      RECT 0.085 2.43 0.465 3.075 ;
      RECT 0.085 2.43 2.595 2.61 ;
      RECT 2.425 1.775 2.595 2.61 ;
      RECT 0.085 1.92 0.455 3.075 ;
      RECT 2.425 1.775 3.01 1.945 ;
      RECT 2.68 1.415 3.01 1.945 ;
      RECT 0.085 0.255 0.26 3.075 ;
      RECT 0.085 0.255 0.425 1.03 ;
      RECT 4.435 2.67 5.495 3 ;
  END
END scs130lp_o21ba_4

MACRO scs130lp_o21ba_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ba_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.115 0.835 1.785 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.115 1.345 1.785 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.82 1.075 3.235 1.745 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.875 2.075 4.205 3.065 ;
        RECT 3.965 0.355 4.205 3.065 ;
        RECT 3.875 0.355 4.205 0.815 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.085 -0.085 3.415 0.815 ;
        RECT 0.66 -0.085 0.99 0.585 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.345 2.785 3.675 3.415 ;
        RECT 1.89 2.785 2.22 3.415 ;
        RECT 0.22 1.965 0.55 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.28 1.965 1.68 2.965 ;
      RECT 1.28 2.435 3.585 2.605 ;
      RECT 3.415 0.995 3.585 2.605 ;
      RECT 1.68 0.265 1.85 2.605 ;
      RECT 3.415 0.995 3.745 1.665 ;
      RECT 1.68 0.265 2.04 0.715 ;
      RECT 2.455 1.925 2.83 2.255 ;
      RECT 2.455 0.355 2.625 2.255 ;
      RECT 2.03 0.905 2.625 1.575 ;
      RECT 2.295 0.355 2.625 1.575 ;
      RECT 0.15 0.765 1.5 0.935 ;
      RECT 1.17 0.265 1.5 0.935 ;
      RECT 0.15 0.265 0.48 0.935 ;
  END
END scs130lp_o21ba_lp

MACRO scs130lp_o21ba_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21ba_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 1.21 3.42 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 2.76 2.49 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.425 1.295 1.75 ;
    END
  END B1N
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.005 0.63 2.86 ;
        RECT 0.155 0.985 0.63 1.195 ;
        RECT 0.155 0.985 0.325 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.965 -0.085 3.175 0.555 ;
        RECT 0.81 0.635 1.02 1.125 ;
        RECT 0.09 0.635 1.02 0.805 ;
        RECT 0.09 -0.085 0.26 0.805 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.995 2.845 3.325 3.415 ;
        RECT 1.835 2.785 2.025 3.415 ;
        RECT 0.885 2.105 1.095 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.555 0.735 3.605 0.905 ;
      RECT 3.395 0.355 3.605 0.905 ;
      RECT 2.555 0.355 2.745 0.905 ;
      RECT 2.205 2.715 2.535 2.925 ;
      RECT 2.205 0.285 2.375 2.925 ;
      RECT 2.045 0.285 2.375 0.495 ;
      RECT 0.44 0.285 2.375 0.455 ;
      RECT 1.335 1.93 1.645 2.94 ;
      RECT 1.475 0.645 1.645 2.94 ;
      RECT 1.475 1.275 2.025 1.445 ;
      RECT 1.855 0.775 2.025 1.445 ;
      RECT 1.255 0.645 1.645 1.195 ;
  END
END scs130lp_o21ba_m

MACRO scs130lp_o21bai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21bai_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.35 1.13 2.795 2.175 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.555 1.13 2.03 1.835 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.035 0.435 2.225 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2905 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.61 2.005 1.905 3.025 ;
        RECT 1.095 2.005 1.905 2.175 ;
        RECT 1.095 0.28 1.465 0.61 ;
        RECT 1.095 0.28 1.385 2.175 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.04 -0.085 2.305 0.61 ;
        RECT 0.585 -0.085 0.915 0.525 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.455 2.345 2.725 3.415 ;
        RECT 1.095 2.345 1.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.635 0.78 2.765 0.95 ;
      RECT 2.475 0.28 2.765 0.95 ;
      RECT 1.635 0.28 1.87 0.95 ;
      RECT 0.615 2.41 0.925 2.74 ;
      RECT 0.675 0.695 0.925 2.74 ;
      RECT 0.155 0.695 0.925 0.865 ;
      RECT 0.155 0.3 0.415 0.865 ;
  END
END scs130lp_o21bai_0

MACRO scs130lp_o21bai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21bai_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.375 2.795 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.58 1.375 2.255 1.75 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.185 0.515 1.89 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7644 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.93 1.925 3.075 ;
        RECT 1.24 1.93 1.925 2.1 ;
        RECT 1.24 0.255 1.41 2.1 ;
        RECT 1.08 0.255 1.41 1.015 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.98 -0.085 2.31 0.865 ;
        RECT 0.525 -0.085 0.855 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.455 1.92 2.785 3.415 ;
        RECT 1.07 2.27 1.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.58 1.035 2.785 1.205 ;
      RECT 2.48 0.255 2.785 1.205 ;
      RECT 1.58 0.255 1.81 1.205 ;
      RECT 0.57 2.06 0.9 2.39 ;
      RECT 0.685 0.845 0.9 2.39 ;
      RECT 0.685 1.185 1.07 1.515 ;
      RECT 0.685 0.845 0.91 1.515 ;
      RECT 0.095 0.845 0.91 1.015 ;
      RECT 0.095 0.385 0.355 1.015 ;
  END
END scs130lp_o21bai_1

MACRO scs130lp_o21bai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21bai_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.515 1.425 3.99 1.645 ;
        RECT 2.015 1.92 3.695 2.12 ;
        RECT 3.515 1.425 3.695 2.12 ;
        RECT 2.015 1.425 2.58 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.8 1.425 3.345 1.75 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.425 1.51 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9408 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 2.29 3.185 2.62 ;
        RECT 1.555 0.595 1.885 1.145 ;
        RECT 1.625 0.595 1.845 2.62 ;
        RECT 1.595 1.815 1.825 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.355 -0.085 3.685 0.915 ;
        RECT 2.435 -0.085 2.765 0.915 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.865 1.815 4.115 3.415 ;
        RECT 1.995 2.79 2.325 3.415 ;
        RECT 0.965 1.815 1.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.065 1.085 4.135 1.255 ;
      RECT 3.855 0.305 4.135 1.255 ;
      RECT 1.125 0.255 1.375 1.185 ;
      RECT 2.935 0.305 3.185 1.255 ;
      RECT 2.065 0.255 2.265 1.255 ;
      RECT 1.125 0.255 2.265 0.425 ;
      RECT 2.495 2.8 3.685 3.075 ;
      RECT 3.355 2.29 3.685 3.075 ;
      RECT 0.46 1.755 0.795 2.21 ;
      RECT 0.595 0.355 0.795 2.21 ;
      RECT 0.595 1.355 1.455 1.605 ;
      RECT 0.595 0.355 0.855 1.605 ;
  END
END scs130lp_o21bai_2

MACRO scs130lp_o21bai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21bai_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.265 1.375 6.615 1.76 ;
        RECT 3.005 1.93 5.435 2.1 ;
        RECT 5.265 1.375 5.435 2.1 ;
        RECT 3.005 1.425 3.335 2.1 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.515 1.425 4.91 1.75 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.415 0.55 1.76 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8816 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.24 2.28 4.79 2.61 ;
        RECT 2.41 2.28 4.79 2.53 ;
        RECT 2.41 0.775 2.725 2.53 ;
        RECT 2.41 0.775 2.6 3.075 ;
        RECT 1.51 1.755 2.725 1.925 ;
        RECT 2.335 0.775 2.725 1.925 ;
        RECT 1.55 0.775 2.725 1.185 ;
        RECT 1.51 1.755 1.74 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.835 -0.085 6.165 0.865 ;
        RECT 4.975 -0.085 5.305 0.845 ;
        RECT 4.115 -0.085 4.445 0.885 ;
        RECT 3.255 -0.085 3.585 0.885 ;
        RECT 0.525 -0.085 0.855 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 6.25 1.93 6.58 3.415 ;
        RECT 5.39 2.63 5.72 3.415 ;
        RECT 2.77 2.7 3.07 3.415 ;
        RECT 1.91 2.105 2.24 3.415 ;
        RECT 0.615 2.27 1.34 3.415 ;
        RECT 1.1 1.825 1.34 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.895 1.055 4.795 1.225 ;
      RECT 6.335 0.255 6.595 1.205 ;
      RECT 4.615 1.035 6.595 1.205 ;
      RECT 3.755 0.255 3.945 1.225 ;
      RECT 2.895 0.255 3.085 1.225 ;
      RECT 4.615 1.015 5.665 1.205 ;
      RECT 5.475 0.255 5.665 1.205 ;
      RECT 4.615 0.255 4.805 1.205 ;
      RECT 1.05 0.255 1.38 0.945 ;
      RECT 1.05 0.255 3.085 0.595 ;
      RECT 5.89 1.93 6.08 3.075 ;
      RECT 3.24 2.79 5.22 3.075 ;
      RECT 4.96 2.27 5.22 3.075 ;
      RECT 4.96 2.27 6.08 2.46 ;
      RECT 5.88 1.93 6.08 2.46 ;
      RECT 0.15 1.93 0.445 3.075 ;
      RECT 0.15 1.93 0.93 2.1 ;
      RECT 0.76 1.075 0.93 2.1 ;
      RECT 0.76 1.325 1.34 1.655 ;
      RECT 0.76 1.355 2.165 1.585 ;
      RECT 0.76 1.325 1.38 1.585 ;
      RECT 0.095 1.075 0.93 1.245 ;
      RECT 0.095 0.255 0.355 1.245 ;
  END
END scs130lp_o21bai_4

MACRO scs130lp_o21bai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21bai_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.27 0.435 2.14 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.27 1.315 2.14 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.25 0.79 2.755 1.12 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3997 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.135 2.31 2.275 2.48 ;
        RECT 1.645 1.55 2.275 2.48 ;
        RECT 1.645 0.595 1.895 2.48 ;
        RECT 1.135 2.31 1.465 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.125 -0.085 2.455 0.61 ;
        RECT 0.635 -0.085 0.965 0.76 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.665 2.66 1.995 3.415 ;
        RECT 0.145 2.31 0.475 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.455 1.33 2.785 3.02 ;
      RECT 2.455 1.33 3.245 1.66 ;
      RECT 3.075 0.295 3.245 1.66 ;
      RECT 2.915 0.295 3.245 0.61 ;
      RECT 0.12 0.93 1.465 1.1 ;
      RECT 1.135 0.605 1.465 1.1 ;
      RECT 0.12 0.605 0.45 1.1 ;
  END
END scs130lp_o21bai_lp

MACRO scs130lp_o21bai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o21bai_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.39 1.21 2.725 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.765 2.12 ;
    END
  END A2
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.505 0.84 0.805 1.51 ;
    END
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.245 2.32 1.765 2.86 ;
        RECT 1.18 2.67 1.415 3 ;
        RECT 1.245 0.5 1.415 3 ;
        RECT 1.205 0.5 1.415 0.83 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 2.065 -0.085 2.275 0.68 ;
        RECT 0.61 -0.085 0.82 0.62 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.97 2.805 2.18 3.415 ;
        RECT 0.66 2.845 0.99 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.635 0.86 2.705 1.03 ;
      RECT 2.495 0.5 2.705 1.03 ;
      RECT 1.635 0.52 1.845 1.03 ;
      RECT 0.15 1.75 0.48 2.925 ;
      RECT 0.895 1.75 1.065 2.42 ;
      RECT 0.15 1.75 1.065 1.92 ;
      RECT 0.15 0.33 0.32 2.925 ;
      RECT 0.15 0.33 0.39 0.66 ;
  END
END scs130lp_o21bai_m

MACRO scs130lp_o221a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221a_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.79 0.78 3.265 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.91 0.765 2.27 1.025 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.535 1.34 2.215 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.535 2.245 2.215 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 1.13 0.865 2.215 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.42 2.63 3.755 2.96 ;
        RECT 3.435 0.28 3.755 2.96 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.935 -0.085 3.265 0.61 ;
        RECT 2.03 -0.085 2.28 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.58 2.725 3.25 3.415 ;
        RECT 0.55 2.725 1.22 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.735 2.385 2.065 3.075 ;
      RECT 0.115 2.385 0.38 3.075 ;
      RECT 0.115 2.385 3.265 2.555 ;
      RECT 2.935 1.93 3.265 2.555 ;
      RECT 0.115 0.575 0.295 3.075 ;
      RECT 0.115 0.575 0.48 0.905 ;
      RECT 1.04 1.195 2.62 1.365 ;
      RECT 2.45 0.28 2.62 1.365 ;
      RECT 1.04 0.61 1.37 1.365 ;
      RECT 2.45 0.28 2.765 0.61 ;
      RECT 1.54 0.255 1.74 0.905 ;
      RECT 0.65 0.255 0.87 0.905 ;
      RECT 0.65 0.255 1.74 0.44 ;
  END
END scs130lp_o221a_0

MACRO scs130lp_o221a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221a_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.955 1.185 3.225 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.185 2.775 1.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.21 1.385 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.195 1.905 1.525 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.345 0.565 1.75 ;
        RECT 0.085 0.755 0.325 2.575 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5817 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.655 2.025 4.235 3.075 ;
        RECT 3.925 0.255 4.235 3.075 ;
        RECT 3.735 1.695 4.235 3.075 ;
        RECT 3.65 0.255 4.235 1.015 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.15 -0.085 3.48 1.015 ;
        RECT 2.29 -0.085 2.62 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.14 2.035 3.47 3.415 ;
        RECT 0.925 2.27 1.255 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.8 1.695 2.63 3.075 ;
      RECT 0.495 1.93 0.755 3.075 ;
      RECT 0.495 1.93 2.63 2.1 ;
      RECT 0.765 1.005 0.935 2.1 ;
      RECT 1.8 1.695 3.565 1.865 ;
      RECT 3.395 1.185 3.565 1.865 ;
      RECT 3.395 1.185 3.755 1.515 ;
      RECT 0.495 1.005 0.935 1.175 ;
      RECT 0.495 0.255 0.73 1.175 ;
      RECT 1.4 0.845 2.98 1.015 ;
      RECT 2.79 0.255 2.98 1.015 ;
      RECT 1.4 0.595 1.6 1.015 ;
      RECT 0.9 0.255 1.23 0.835 ;
      RECT 1.77 0.255 2.1 0.675 ;
      RECT 0.9 0.255 2.1 0.425 ;
  END
END scs130lp_o221a_1

MACRO scs130lp_o221a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221a_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.345 2.955 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.335 2.375 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.885 1.345 1.295 1.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.335 1.805 1.75 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.375 1.76 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.48 1.815 4.22 1.985 ;
        RECT 3.77 1.065 4.22 1.985 ;
        RECT 3.425 1.065 4.22 1.235 ;
        RECT 3.425 0.255 3.685 1.235 ;
        RECT 3.48 1.815 3.67 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.855 -0.085 4.155 0.895 ;
        RECT 3.01 -0.085 3.255 1.095 ;
        RECT 2.03 -0.085 2.36 0.825 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.84 2.165 4.17 3.415 ;
        RECT 2.64 2.27 3.31 3.415 ;
        RECT 0.665 2.27 0.995 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.51 1.93 2.195 3.075 ;
      RECT 0.18 1.93 0.495 3.075 ;
      RECT 0.18 1.93 3.295 2.1 ;
      RECT 3.125 1.405 3.295 2.1 ;
      RECT 0.545 0.86 0.715 2.1 ;
      RECT 3.125 1.405 3.6 1.645 ;
      RECT 0.14 0.86 0.715 1.03 ;
      RECT 0.14 0.315 0.4 1.03 ;
      RECT 1.07 0.995 2.84 1.165 ;
      RECT 2.53 0.255 2.84 1.165 ;
      RECT 1.07 0.595 1.4 1.165 ;
      RECT 1.57 0.255 1.84 0.825 ;
      RECT 0.57 0.255 0.9 0.69 ;
      RECT 0.57 0.255 1.84 0.425 ;
  END
END scs130lp_o221a_2

MACRO scs130lp_o221a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221a_4 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.465 1.075 5.03 1.515 ;
        RECT 3.37 1.075 5.03 1.245 ;
        RECT 3.37 1.075 3.69 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.86 1.425 4.295 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.075 3.155 1.605 ;
        RECT 1.595 1.075 3.155 1.245 ;
        RECT 1.035 1.21 1.82 1.605 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 1.425 2.735 1.76 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.35 0.435 1.785 ;
        RECT 0.085 1.21 0.35 1.785 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.54 1.755 7.115 1.925 ;
        RECT 6.865 1.045 7.115 1.925 ;
        RECT 5.465 1.045 7.115 1.215 ;
        RECT 6.4 1.755 6.59 3.075 ;
        RECT 6.365 0.255 6.555 1.215 ;
        RECT 5.54 1.755 5.73 3.075 ;
        RECT 5.465 0.255 5.695 1.215 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 6.725 -0.085 7.055 0.875 ;
        RECT 5.865 -0.085 6.195 0.865 ;
        RECT 5.035 -0.085 5.295 0.905 ;
        RECT 4.105 -0.085 4.435 0.54 ;
        RECT 3.245 -0.085 3.575 0.54 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 6.76 2.105 7.09 3.415 ;
        RECT 5.9 2.105 6.23 3.415 ;
        RECT 4.97 2.27 5.3 3.415 ;
        RECT 2.725 2.27 3.505 3.415 ;
        RECT 0.985 2.27 1.315 3.415 ;
        RECT 0.105 1.955 0.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.605 0.595 0.815 3.075 ;
      RECT 4.035 1.93 4.365 2.735 ;
      RECT 1.865 1.93 2.195 2.735 ;
      RECT 0.605 1.93 5.37 2.1 ;
      RECT 5.2 1.385 5.37 2.1 ;
      RECT 0.605 0.595 0.865 2.1 ;
      RECT 5.2 1.385 6.695 1.585 ;
      RECT 0.535 0.595 0.865 1.145 ;
      RECT 1.435 0.725 4.865 0.905 ;
      RECT 3.135 0.71 4.865 0.905 ;
      RECT 1.435 0.71 2.645 0.905 ;
      RECT 3.675 2.905 4.795 3.075 ;
      RECT 4.535 2.28 4.795 3.075 ;
      RECT 3.675 2.27 3.865 3.075 ;
      RECT 0.105 0.255 0.365 1.04 ;
      RECT 1.035 0.255 1.265 0.975 ;
      RECT 2.725 0.255 3.055 0.555 ;
      RECT 1.035 0.255 3.055 0.54 ;
      RECT 0.105 0.255 3.055 0.425 ;
      RECT 1.485 2.905 2.555 3.075 ;
      RECT 2.365 2.27 2.555 3.075 ;
      RECT 1.485 2.27 1.695 3.075 ;
  END
END scs130lp_o221a_4

MACRO scs130lp_o221a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221a_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.02 1.12 1.35 1.79 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.12 1.87 1.79 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.33 3.33 1.78 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.04 1.395 2.765 1.78 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.5 1.33 3.895 1.79 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 2.075 0.49 3.065 ;
        RECT 0.1 0.265 0.445 1.04 ;
        RECT 0.1 0.265 0.27 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 1.845 -0.085 2.175 0.365 ;
        RECT 0.905 -0.085 1.155 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 2.875 2.32 3.205 3.415 ;
        RECT 0.69 2.32 1.02 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.405 1.97 4.235 3.065 ;
      RECT 4.065 0.685 4.235 3.065 ;
      RECT 1.815 1.97 2.145 3.065 ;
      RECT 0.67 1.97 4.235 2.14 ;
      RECT 0.67 1.225 0.84 2.14 ;
      RECT 0.45 1.225 0.84 1.895 ;
      RECT 3.865 0.685 4.235 1.015 ;
      RECT 2.425 0.99 3.695 1.16 ;
      RECT 3.445 0.685 3.695 1.16 ;
      RECT 2.425 0.895 2.755 1.16 ;
      RECT 2.935 0.545 3.265 0.82 ;
      RECT 1.335 0.545 3.265 0.715 ;
      RECT 1.335 0.265 1.665 0.715 ;
  END
END scs130lp_o221a_lp

MACRO scs130lp_o221a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221a_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.3 1.09 2.775 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.845 2.01 2.515 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.925 0.925 2.12 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.815 1.415 2.145 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 0.39 0.855 0.72 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.95 2.655 3.26 2.985 ;
        RECT 3.09 0.345 3.26 2.985 ;
        RECT 2.995 0.345 3.26 1.75 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.565 -0.085 2.775 0.545 ;
        RECT 1.625 -0.085 1.955 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.54 2.785 2.73 3.415 ;
        RECT 0.65 2.845 0.98 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.245 2.695 2.36 3.025 ;
      RECT 2.19 1.97 2.36 3.025 ;
      RECT 0.14 2.495 0.47 2.925 ;
      RECT 1.245 2.495 1.415 3.025 ;
      RECT 0.14 2.495 1.415 2.665 ;
      RECT 0.14 1.005 0.365 2.925 ;
      RECT 2.19 1.97 2.91 2.3 ;
      RECT 1.05 0.665 1.38 1.145 ;
      RECT 1.05 0.665 2.345 0.835 ;
      RECT 2.135 0.345 2.345 0.835 ;
      RECT 0.585 1.325 1.845 1.495 ;
      RECT 1.635 1.035 1.845 1.495 ;
      RECT 0.585 1.005 0.795 1.495 ;
  END
END scs130lp_o221a_m

MACRO scs130lp_o221ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221ai_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.46 1.42 3.27 1.755 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.46 1.31 2.28 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.21 1.29 1.76 ;
        RECT 0.545 1.21 1.29 1.41 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.955 1.93 3.275 2.945 ;
        RECT 1.105 1.93 3.275 2.14 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.92 0.585 2.15 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5305 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 2.32 1.795 2.99 ;
        RECT 0.185 2.32 1.795 2.49 ;
        RECT 0.765 1.58 0.935 2.49 ;
        RECT 0.095 1.58 0.935 1.75 ;
        RECT 0.185 2.32 0.445 3 ;
        RECT 0.095 0.28 0.365 1.75 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.465 -0.085 2.135 0.36 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.365 2.33 2.695 3.415 ;
        RECT 0.615 2.66 0.945 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.465 0.875 3.075 1.045 ;
      RECT 2.77 0.28 3.075 1.045 ;
      RECT 0.545 0.87 1.635 1.04 ;
      RECT 0.545 0.28 0.715 1.04 ;
      RECT 0.545 0.28 0.835 0.615 ;
      RECT 1.005 0.53 2.6 0.7 ;
      RECT 2.315 0.28 2.6 0.7 ;
      RECT 1.005 0.28 1.285 0.7 ;
  END
END scs130lp_o221ai_0

MACRO scs130lp_o221ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221ai_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.345 3.275 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.49 1.345 2.735 2.96 ;
        RECT 2.27 1.345 2.735 1.675 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.345 1.375 1.78 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.345 2.06 1.775 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.345 0.455 1.76 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2747 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 1.95 2.32 3.075 ;
        RECT 0.295 1.95 2.32 2.12 ;
        RECT 0.295 1.93 0.885 2.12 ;
        RECT 0.625 1.005 0.885 2.12 ;
        RECT 0.115 1.005 0.885 1.175 ;
        RECT 0.295 1.93 0.555 3.075 ;
        RECT 0.115 0.255 0.375 1.175 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.495 -0.085 2.825 0.835 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.935 1.92 3.265 3.415 ;
        RECT 0.725 2.29 1.395 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.065 1.005 3.265 1.175 ;
      RECT 2.995 0.255 3.265 1.175 ;
      RECT 1.065 0.995 2.325 1.175 ;
      RECT 2.05 0.255 2.325 1.175 ;
      RECT 1.065 0.595 1.38 1.175 ;
      RECT 0.545 0.255 0.875 0.835 ;
      RECT 1.55 0.255 1.88 0.815 ;
      RECT 0.545 0.255 1.88 0.425 ;
  END
END scs130lp_o221ai_1

MACRO scs130lp_o221ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221ai_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.68 1.695 5.67 1.875 ;
        RECT 5.345 1.21 5.67 1.875 ;
        RECT 3.68 1.345 4.015 1.875 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.22 1.21 5.175 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.505 1.705 3.47 1.875 ;
        RECT 3.14 1.345 3.47 1.875 ;
        RECT 1.505 1.425 2.315 1.875 ;
        RECT 1.35 1.425 2.315 1.675 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.485 1.21 2.835 1.535 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 1.21 0.355 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2936 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.455 2.045 4.785 2.725 ;
        RECT 0.535 2.045 4.785 2.215 ;
        RECT 2.415 2.045 2.745 2.735 ;
        RECT 0.535 1.845 1.335 2.215 ;
        RECT 0.535 1.815 1.18 2.215 ;
        RECT 0.535 0.595 0.865 2.215 ;
        RECT 0.535 0.595 0.795 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.795 -0.085 5.125 0.7 ;
        RECT 3.895 -0.085 4.225 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.315 2.045 5.645 3.415 ;
        RECT 3.395 2.385 3.725 3.415 ;
        RECT 0.965 2.385 1.815 3.415 ;
        RECT 0.105 1.92 0.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.515 0.87 5.575 1.04 ;
      RECT 5.295 0.305 5.575 1.04 ;
      RECT 1.485 0.255 1.815 0.915 ;
      RECT 4.395 0.305 4.625 1.04 ;
      RECT 3.515 0.255 3.715 1.04 ;
      RECT 2.485 0.255 2.695 0.7 ;
      RECT 1.485 0.255 3.715 0.425 ;
      RECT 4.025 2.895 5.145 3.075 ;
      RECT 4.955 2.045 5.145 3.075 ;
      RECT 4.025 2.385 4.285 3.075 ;
      RECT 1.045 1.085 2.315 1.255 ;
      RECT 1.985 0.595 2.315 1.255 ;
      RECT 3.005 0.595 3.345 1.145 ;
      RECT 1.045 0.255 1.235 1.255 ;
      RECT 1.985 0.87 3.345 1.04 ;
      RECT 2.865 0.595 3.345 1.04 ;
      RECT 0.105 0.255 0.365 1.04 ;
      RECT 0.105 0.255 1.235 0.425 ;
      RECT 1.985 2.905 3.175 3.075 ;
      RECT 2.915 2.385 3.175 3.075 ;
      RECT 1.985 2.385 2.245 3.075 ;
  END
END scs130lp_o221ai_2

MACRO scs130lp_o221ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221ai_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.385 1.21 9.99 1.52 ;
        RECT 6.405 1.075 8.59 1.245 ;
        RECT 6.405 1.075 6.655 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.825 1.425 8.215 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.81 1.615 6.145 1.785 ;
        RECT 5.815 1.295 6.145 1.785 ;
        RECT 2.81 1.4 3.82 1.785 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.225 1.195 5.645 1.445 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.425 2.29 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.6544 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.85 1.95 8.18 2.735 ;
        RECT 6.395 1.95 8.18 2.12 ;
        RECT 6.99 1.95 7.32 2.735 ;
        RECT 4.225 1.955 7.32 2.135 ;
        RECT 5.085 1.955 5.415 2.735 ;
        RECT 4.225 1.955 4.555 2.735 ;
        RECT 2.145 1.955 7.32 2.125 ;
        RECT 1.285 1.92 2.64 2.09 ;
        RECT 2.46 1.085 2.64 2.125 ;
        RECT 0.535 1.085 2.64 1.255 ;
        RECT 2.145 1.92 2.335 3.075 ;
        RECT 1.535 0.595 1.865 1.255 ;
        RECT 1.285 1.92 1.465 3.075 ;
        RECT 0.535 0.595 0.865 1.255 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.14 -0.085 9.47 0.7 ;
        RECT 8.28 -0.085 8.61 0.565 ;
        RECT 7.42 -0.085 7.75 0.565 ;
        RECT 6.56 -0.085 6.89 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.64 1.815 9.935 3.415 ;
        RECT 8.745 2.03 9.075 3.415 ;
        RECT 6.05 2.305 6.38 3.415 ;
        RECT 3.365 2.635 3.695 3.415 ;
        RECT 2.505 2.295 2.835 3.415 ;
        RECT 1.645 2.26 1.975 3.415 ;
        RECT 0.785 1.92 1.115 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.76 0.87 9.9 1.04 ;
      RECT 9.64 0.255 9.9 1.04 ;
      RECT 6.06 0.255 6.29 0.945 ;
      RECT 6.06 0.735 8.97 0.905 ;
      RECT 3.365 0.255 3.695 0.835 ;
      RECT 8.78 0.255 8.97 1.04 ;
      RECT 7.92 0.255 8.11 0.905 ;
      RECT 7.06 0.255 7.25 0.905 ;
      RECT 6.06 0.255 6.39 0.905 ;
      RECT 4.285 0.255 5.355 0.605 ;
      RECT 2.505 0.255 3.695 0.485 ;
      RECT 2.505 0.255 6.39 0.445 ;
      RECT 9.245 1.69 9.47 3.075 ;
      RECT 6.56 2.905 8.575 3.075 ;
      RECT 8.385 1.69 8.575 3.075 ;
      RECT 7.49 2.29 7.68 3.075 ;
      RECT 6.56 2.305 6.82 3.075 ;
      RECT 8.385 1.69 9.47 1.86 ;
      RECT 2.81 1.005 4.045 1.23 ;
      RECT 0.105 0.255 0.365 1.185 ;
      RECT 5.515 0.665 5.845 1.025 ;
      RECT 3.865 0.775 5.845 1.025 ;
      RECT 2.81 0.655 3.195 1.23 ;
      RECT 2.035 0.655 3.195 0.915 ;
      RECT 1.035 0.255 1.365 0.895 ;
      RECT 3.865 0.615 4.115 1.025 ;
      RECT 2.035 0.255 2.315 0.915 ;
      RECT 0.105 0.255 2.315 0.425 ;
      RECT 3.865 2.905 5.845 3.075 ;
      RECT 5.585 2.305 5.845 3.075 ;
      RECT 3.005 2.295 3.195 3.075 ;
      RECT 4.725 2.315 4.915 3.075 ;
      RECT 3.865 2.295 4.055 3.075 ;
      RECT 3.005 2.295 4.055 2.465 ;
  END
END scs130lp_o221ai_4

MACRO scs130lp_o221ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221ai_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 0.915 3.265 1.585 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.02 1.035 2.755 1.41 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.405 1.18 1.795 1.85 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.765 3.835 1.935 ;
        RECT 3.485 0.895 3.835 1.935 ;
        RECT 1.975 1.605 2.305 1.935 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 1.05 0.875 1.72 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7247 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.2 2.465 2.53 3.065 ;
        RECT 0.125 2.465 2.53 2.635 ;
        RECT 0.125 1.92 0.875 3.065 ;
        RECT 0.125 0.265 0.875 0.715 ;
        RECT 0.125 0.265 0.295 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 2.075 -0.085 2.405 0.505 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.26 2.465 3.59 3.415 ;
        RECT 1.075 2.815 1.405 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.055 2.115 4.185 2.285 ;
      RECT 4.015 0.265 4.185 2.285 ;
      RECT 1.055 0.265 1.225 2.285 ;
      RECT 1.055 0.265 1.385 0.895 ;
      RECT 3.71 0.265 4.185 0.715 ;
      RECT 1.565 0.685 2.755 0.855 ;
      RECT 3.2 0.265 3.53 0.715 ;
      RECT 2.585 0.545 3.53 0.715 ;
      RECT 1.565 0.265 1.895 0.855 ;
  END
END scs130lp_o221ai_lp

MACRO scs130lp_o221ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o221ai_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.535 1.885 3.205 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 0.995 1.795 1.505 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 1.21 1.285 1.405 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.84 2.905 1.355 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.505 1.95 0.835 2.12 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.44125 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.715 2.3 1.925 2.63 ;
        RECT 0.155 2.3 1.925 2.47 ;
        RECT 0.155 0.345 0.555 0.675 ;
        RECT 0.155 2.3 0.49 2.86 ;
        RECT 0.155 0.345 0.325 2.86 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.61 -0.085 1.94 0.465 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.54 2.485 2.87 3.415 ;
        RECT 0.71 2.65 1.04 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.015 1.685 2.145 1.855 ;
      RECT 0.545 1.585 1.185 1.755 ;
      RECT 3.085 0.33 3.255 1.705 ;
      RECT 1.975 1.535 3.255 1.705 ;
      RECT 0.545 0.86 0.715 1.755 ;
      RECT 0.545 0.86 0.985 1.03 ;
      RECT 0.775 0.345 0.985 1.03 ;
      RECT 2.65 0.33 3.255 0.66 ;
      RECT 1.22 0.645 2.375 0.815 ;
      RECT 2.205 0.33 2.43 0.66 ;
      RECT 1.22 0.345 1.43 0.815 ;
  END
END scs130lp_o221ai_m

MACRO scs130lp_o22a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22a_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 2.095 3.37 2.265 ;
        RECT 3.06 1.935 3.37 2.265 ;
        RECT 1.515 1.215 1.685 2.265 ;
        RECT 0.99 1.215 1.685 1.395 ;
        RECT 0.995 0.265 1.325 0.435 ;
        RECT 0.99 1.17 1.295 1.395 ;
        RECT 1.115 0.265 1.295 1.395 ;
        RECT 0.995 0.265 1.295 0.5 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.245 1.115 3.755 1.415 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.565 1.345 2.235 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.955 1.385 2.735 1.925 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.605 0.465 0.935 ;
        RECT 0.085 2.425 0.425 3.075 ;
        RECT 0.085 0.605 0.325 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.875 -0.085 3.205 0.865 ;
        RECT 0.645 0.67 0.945 1 ;
        RECT 0.645 -0.085 0.825 1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.185 2.775 3.515 3.415 ;
        RECT 0.595 2.775 1.735 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.225 2.435 2.555 3.075 ;
      RECT 0.595 2.435 3.745 2.605 ;
      RECT 3.54 1.585 3.745 2.605 ;
      RECT 0.595 2.065 0.765 2.605 ;
      RECT 0.495 1.565 0.665 2.235 ;
      RECT 2.905 1.585 3.745 1.755 ;
      RECT 2.905 1.035 3.075 1.755 ;
      RECT 1.855 1.035 3.075 1.205 ;
      RECT 1.855 0.785 2.185 1.205 ;
      RECT 1.465 0.615 1.685 1 ;
      RECT 2.365 0.445 2.695 0.865 ;
      RECT 1.495 0.445 2.695 0.615 ;
  END
END scs130lp_o22a_0

MACRO scs130lp_o22a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22a_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.375 3.715 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.425 3.205 2.86 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.41 1.425 1.765 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 1.425 2.31 1.75 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.67 1.815 0.88 2.825 ;
        RECT 0.155 1.815 0.88 1.985 ;
        RECT 0.155 0.425 0.365 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.7 -0.085 3.03 0.825 ;
        RECT 0.585 -0.085 0.795 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.385 2.105 3.595 3.415 ;
        RECT 1.1 2.445 1.31 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.225 1.005 3.54 1.175 ;
      RECT 3.33 0.425 3.54 1.175 ;
      RECT 2.225 0.345 2.435 1.175 ;
      RECT 1.285 0.345 1.615 0.895 ;
      RECT 1.285 0.345 2.435 0.515 ;
      RECT 2.165 1.93 2.375 2.94 ;
      RECT 1.06 1.93 2.375 2.1 ;
      RECT 1.06 1.075 1.23 2.1 ;
      RECT 0.55 1.075 0.88 1.435 ;
      RECT 0.55 1.075 2.005 1.245 ;
      RECT 1.795 0.765 2.005 1.245 ;
  END
END scs130lp_o22a_1

MACRO scs130lp_o22a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22a_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.375 3.755 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.76 1.345 3.205 2.94 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.48 1.425 1.895 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.425 2.47 1.75 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.62 1.075 0.88 3.075 ;
        RECT 0.535 0.255 0.775 1.825 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.875 -0.085 3.205 0.825 ;
        RECT 0.955 -0.085 1.285 0.905 ;
        RECT 0.095 -0.085 0.365 1.105 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.375 1.92 3.69 3.415 ;
        RECT 1.06 2.27 1.805 3.415 ;
        RECT 0.2 1.995 0.45 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.375 0.995 3.69 1.165 ;
      RECT 3.375 0.255 3.69 1.165 ;
      RECT 2.375 0.255 2.705 1.165 ;
      RECT 1.475 0.255 1.805 0.895 ;
      RECT 1.475 0.255 2.705 0.425 ;
      RECT 2.245 1.93 2.59 3.075 ;
      RECT 1.05 1.93 2.59 2.1 ;
      RECT 1.05 1.075 1.31 2.1 ;
      RECT 1.05 1.075 2.205 1.245 ;
      RECT 1.975 0.595 2.205 1.245 ;
  END
END scs130lp_o22a_2

MACRO scs130lp_o22a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22a_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.85 1.185 6.625 1.77 ;
        RECT 4.65 1.075 6.055 1.245 ;
        RECT 4.65 1.075 4.98 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.19 1.425 5.68 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.11 1.075 4.44 1.515 ;
        RECT 3.035 1.075 4.44 1.245 ;
        RECT 2.86 1.195 3.285 1.525 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.455 1.415 3.9 1.76 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.15 1.755 2.34 3.075 ;
        RECT 0.085 1.755 2.34 1.925 ;
        RECT 0.085 1.055 1.715 1.225 ;
        RECT 1.485 0.255 1.715 1.225 ;
        RECT 1.29 1.755 1.48 3.075 ;
        RECT 0.625 0.255 0.815 1.225 ;
        RECT 0.085 1.055 0.505 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.745 -0.085 6.075 0.565 ;
        RECT 4.845 -0.085 5.175 0.565 ;
        RECT 1.885 -0.085 2.125 1.105 ;
        RECT 0.985 -0.085 1.315 0.885 ;
        RECT 0.125 -0.085 0.455 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 6.175 1.94 6.505 3.415 ;
        RECT 4.38 2.27 4.71 3.415 ;
        RECT 2.545 2.27 2.875 3.415 ;
        RECT 1.65 2.105 1.98 3.415 ;
        RECT 0.79 2.095 1.12 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.225 0.735 6.505 1.015 ;
      RECT 6.245 0.255 6.505 1.015 ;
      RECT 2.635 0.685 2.865 1.015 ;
      RECT 2.635 0.735 6.505 0.905 ;
      RECT 5.345 0.255 5.575 0.905 ;
      RECT 2.635 0.685 4.675 0.905 ;
      RECT 4.385 0.255 4.675 0.905 ;
      RECT 4.885 2.905 6.005 3.075 ;
      RECT 5.815 1.94 6.005 3.075 ;
      RECT 4.885 2.27 5.145 3.075 ;
      RECT 5.315 1.93 5.645 2.735 ;
      RECT 3.445 1.93 3.775 2.735 ;
      RECT 2.51 1.93 5.645 2.1 ;
      RECT 2.51 1.405 2.68 2.1 ;
      RECT 0.775 1.405 2.68 1.575 ;
      RECT 2.295 0.255 2.465 1.575 ;
      RECT 2.295 0.255 4.205 0.515 ;
      RECT 3.045 2.905 4.205 3.075 ;
      RECT 3.945 2.27 4.205 3.075 ;
      RECT 3.045 2.27 3.275 3.075 ;
  END
END scs130lp_o22a_4

MACRO scs130lp_o22a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22a_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.11 1.585 0.615 2.14 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.825 1.585 1.33 2.14 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.115 1.45 2.755 1.78 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 0.325 2.275 0.67 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.285 2.075 3.725 3.065 ;
        RECT 3.485 0.265 3.725 3.065 ;
        RECT 3.395 0.265 3.725 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.605 -0.085 2.935 0.615 ;
        RECT 0.575 -0.085 0.905 1.075 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.22 2.31 2.55 3.415 ;
        RECT 0.115 2.31 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.135 2.31 1.465 3.065 ;
      RECT 1.135 2.31 1.855 2.48 ;
      RECT 1.685 1.2 1.855 2.48 ;
      RECT 1.685 1.96 3.105 2.13 ;
      RECT 2.935 0.855 3.105 2.13 ;
      RECT 1.685 1.2 1.935 2.13 ;
      RECT 2.935 0.855 3.265 1.525 ;
      RECT 0.13 1.245 1.505 1.415 ;
      RECT 1.095 0.85 1.505 1.415 ;
      RECT 2.115 0.85 2.445 1.27 ;
      RECT 0.13 0.85 0.405 1.415 ;
      RECT 1.095 0.85 2.445 1.02 ;
  END
END scs130lp_o22a_lp

MACRO scs130lp_o22a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22a_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.885 1.495 3.205 2.49 ;
        RECT 1.005 1.495 3.205 1.665 ;
        RECT 1.005 1.165 1.335 1.675 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.485 0.84 3.205 1.185 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.95 1.285 2.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.845 2.245 2.355 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.14 0.445 0.47 0.635 ;
        RECT 0.14 0.445 0.365 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.69 -0.085 3.02 0.655 ;
        RECT 0.65 -0.085 0.98 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.93 2.845 3.26 3.415 ;
        RECT 0.565 2.885 0.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.18 0.265 2.51 0.655 ;
      RECT 1.16 0.265 1.49 0.635 ;
      RECT 1.16 0.265 2.51 0.435 ;
      RECT 2.09 2.535 2.3 2.985 ;
      RECT 0.545 2.535 2.3 2.705 ;
      RECT 0.545 0.815 0.715 2.705 ;
      RECT 0.545 0.815 2 0.985 ;
      RECT 1.67 0.615 2 0.985 ;
  END
END scs130lp_o22a_m

MACRO scs130lp_o22ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22ai_0 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 1.21 2.315 2.205 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.21 1.83 2.13 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.385 2.12 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 1.21 1.295 2.12 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3283 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.08 2.3 1.765 3.065 ;
        RECT 0.555 2.3 1.765 2.49 ;
        RECT 0.625 0.595 0.955 1.005 ;
        RECT 0.555 0.835 0.725 2.49 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.525 -0.085 1.855 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.935 2.395 2.23 3.415 ;
        RECT 0.125 2.66 0.59 3.415 ;
        RECT 0.125 2.395 0.385 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.135 0.87 2.305 1.04 ;
      RECT 2.025 0.47 2.305 1.04 ;
      RECT 1.135 0.255 1.355 1.04 ;
      RECT 0.115 0.255 0.445 0.67 ;
      RECT 0.115 0.255 1.355 0.425 ;
  END
END scs130lp_o22ai_0

MACRO scs130lp_o22ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22ai_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.795 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.455 1.21 1.765 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.355 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.865 1.345 1.285 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0479 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.525 1.93 1.6 3.075 ;
        RECT 0.525 0.595 0.855 1.175 ;
        RECT 0.525 0.595 0.695 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.45 -0.085 2.12 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.04 1.92 2.37 3.415 ;
        RECT 0.095 1.92 0.355 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.025 0.87 2.55 1.04 ;
      RECT 2.29 0.325 2.55 1.04 ;
      RECT 0.095 0.255 0.355 1.04 ;
      RECT 1.025 0.255 1.28 1.04 ;
      RECT 0.095 0.255 1.28 0.425 ;
  END
END scs130lp_o22ai_1

MACRO scs130lp_o22ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22ai_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.94 1.21 4.715 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.45 1.21 3.77 1.525 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.355 0.935 1.605 ;
        RECT 0.155 1.21 0.435 1.605 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 1.21 1.83 1.525 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.845 1.695 3.175 2.735 ;
        RECT 1.465 1.695 3.175 1.865 ;
        RECT 2 0.82 2.255 1.865 ;
        RECT 0.605 0.82 2.255 1.03 ;
        RECT 1.465 1.695 1.795 2.735 ;
        RECT 0.605 0.595 0.935 1.185 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.635 -0.085 3.965 0.7 ;
        RECT 2.775 -0.085 3.105 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.705 2.035 4.035 3.415 ;
        RECT 0.605 2.115 0.935 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.205 1.695 4.465 3.075 ;
      RECT 2.415 2.905 3.535 3.075 ;
      RECT 3.345 1.695 3.535 3.075 ;
      RECT 2.415 2.035 2.675 3.075 ;
      RECT 3.345 1.695 4.465 1.865 ;
      RECT 2.425 0.87 4.395 1.04 ;
      RECT 4.135 0.315 4.395 1.04 ;
      RECT 0.175 0.255 0.435 1.04 ;
      RECT 3.285 0.315 3.465 1.04 ;
      RECT 2.425 0.255 2.605 1.04 ;
      RECT 1.105 0.255 2.605 0.65 ;
      RECT 0.175 0.255 2.605 0.425 ;
      RECT 1.105 2.905 2.225 3.075 ;
      RECT 1.965 2.035 2.225 3.075 ;
      RECT 0.175 1.775 0.435 3.075 ;
      RECT 1.105 1.775 1.295 3.075 ;
      RECT 0.175 1.775 1.295 1.945 ;
  END
END scs130lp_o22ai_2

MACRO scs130lp_o22ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22ai_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.345 3.715 1.525 ;
        RECT 1.025 1.95 3.555 2.12 ;
        RECT 3.385 1.345 3.555 2.12 ;
        RECT 1.025 1.345 1.455 2.12 ;
        RECT 0.105 1.345 1.455 1.63 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.81 1.345 3.205 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.93 1.005 7.195 1.515 ;
        RECT 4.885 1.005 7.195 1.175 ;
        RECT 3.955 1.355 5.125 1.535 ;
        RECT 4.885 1.005 5.125 1.535 ;
        RECT 3.995 1.21 5.125 1.535 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.305 1.345 6.655 1.535 ;
        RECT 5.81 1.345 6.12 1.76 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.29 1.705 7.535 1.875 ;
        RECT 7.365 0.645 7.535 1.875 ;
        RECT 3.985 0.645 7.535 0.835 ;
        RECT 6.23 1.93 6.56 2.735 ;
        RECT 6.29 1.705 6.56 2.735 ;
        RECT 5.37 1.93 6.56 2.1 ;
        RECT 5.37 1.93 5.7 2.735 ;
        RECT 5.37 1.705 5.64 2.735 ;
        RECT 3.79 1.705 5.64 1.875 ;
        RECT 3.985 0.645 4.715 1.04 ;
        RECT 1.92 2.29 3.96 2.47 ;
        RECT 3.79 1.705 3.96 2.47 ;
        RECT 1.92 2.29 3.05 2.62 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 3.135 -0.085 3.465 0.825 ;
        RECT 2.275 -0.085 2.605 0.825 ;
        RECT 1.415 -0.085 1.745 0.825 ;
        RECT 0.555 -0.085 0.885 0.825 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 7.09 2.105 7.42 3.415 ;
        RECT 4.51 2.395 4.84 3.415 ;
        RECT 3.65 2.64 3.96 3.415 ;
        RECT 1 2.63 1.33 3.415 ;
        RECT 0.14 1.815 0.43 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.125 1.005 3.815 1.175 ;
      RECT 3.635 0.255 3.815 1.175 ;
      RECT 2.775 0.255 2.965 1.175 ;
      RECT 1.915 0.255 2.105 1.175 ;
      RECT 1.055 0.255 1.245 1.175 ;
      RECT 0.125 0.255 0.385 1.175 ;
      RECT 3.635 0.255 7.39 0.475 ;
      RECT 5.01 2.905 6.92 3.075 ;
      RECT 6.73 2.045 6.92 3.075 ;
      RECT 4.13 2.045 4.34 3.075 ;
      RECT 5.87 2.27 6.06 3.075 ;
      RECT 5.01 2.045 5.2 3.075 ;
      RECT 4.13 2.045 5.2 2.225 ;
      RECT 1.5 2.79 3.48 3.075 ;
      RECT 0.6 1.815 0.83 3.075 ;
      RECT 1.5 2.29 1.7 3.075 ;
      RECT 0.6 2.29 1.7 2.46 ;
      RECT 0.6 1.815 0.855 2.46 ;
  END
END scs130lp_o22ai_4

MACRO scs130lp_o22ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22ai_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 1.035 2.845 1.705 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 1.035 2.275 1.705 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.515 1.45 0.845 1.78 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.45 1.415 1.78 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 2.235 1.64 3.065 ;
        RECT 1.085 1.96 1.315 3.065 ;
        RECT 0.165 1.1 1.17 1.27 ;
        RECT 0.84 0.615 1.17 1.27 ;
        RECT 0.165 1.96 1.315 2.13 ;
        RECT 0.165 1.1 0.335 2.13 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.945 -0.085 2.275 0.855 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.74 2.235 3.07 3.415 ;
        RECT 0.29 2.31 0.62 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.595 1.885 3.195 2.055 ;
      RECT 3.025 0.485 3.195 2.055 ;
      RECT 1.595 0.265 1.765 2.055 ;
      RECT 1.35 0.265 1.765 0.945 ;
      RECT 0.33 0.265 0.66 0.92 ;
      RECT 2.64 0.485 3.195 0.855 ;
      RECT 0.33 0.265 1.765 0.435 ;
  END
END scs130lp_o22ai_lp

MACRO scs130lp_o22ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o22ai_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.41 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.84 2.12 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.86 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.1 1.21 1.285 2.12 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2352 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 2.715 1.655 2.925 ;
        RECT 1.115 2.32 1.285 2.925 ;
        RECT 0.895 0.62 1.225 1.01 ;
        RECT 0.75 2.32 1.285 2.49 ;
        RECT 0.75 0.84 0.92 2.49 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.855 -0.085 2.185 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.115 2.845 2.445 3.415 ;
        RECT 0.535 2.845 0.865 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.465 0.84 2.555 1.01 ;
      RECT 2.365 0.52 2.555 1.01 ;
      RECT 1.465 0.27 1.675 1.01 ;
      RECT 0.385 0.27 0.715 0.66 ;
      RECT 0.385 0.27 1.675 0.44 ;
  END
END scs130lp_o22ai_m

MACRO scs130lp_o2bb2a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2a_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.885 1.55 1.295 2.13 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1 1.015 1.61 1.38 ;
        RECT 1 0.86 1.35 1.38 ;
        RECT 1.105 0.395 1.35 1.38 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.2 1.155 3.755 2.215 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.155 2.99 1.825 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 0.38 0.505 0.71 ;
        RECT 0.095 2.395 0.355 3.065 ;
        RECT 0.095 0.38 0.325 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3 -0.085 3.26 0.61 ;
        RECT 0.675 -0.085 0.935 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.325 2.46 3.655 3.415 ;
        RECT 2.145 2.515 2.405 3.415 ;
        RECT 0.525 2.64 0.835 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.545 0.78 3.725 0.95 ;
      RECT 3.43 0.28 3.725 0.95 ;
      RECT 2.545 0.28 2.83 0.95 ;
      RECT 1.005 2.905 1.975 3.075 ;
      RECT 1.805 2.175 1.975 3.075 ;
      RECT 1.005 2.3 1.175 3.075 ;
      RECT 2.575 2.175 2.865 2.79 ;
      RECT 0.545 2.3 1.175 2.47 ;
      RECT 1.805 2.175 2.865 2.345 ;
      RECT 0.545 0.88 0.715 2.47 ;
      RECT 2.205 0.28 2.375 2.345 ;
      RECT 0.495 0.88 0.715 1.55 ;
      RECT 2.13 0.28 2.375 0.675 ;
      RECT 1.345 2.405 1.635 2.735 ;
      RECT 1.465 1.745 1.635 2.735 ;
      RECT 1.465 1.745 2.035 1.915 ;
      RECT 1.79 1.585 2.035 1.915 ;
      RECT 1.79 0.395 1.96 1.915 ;
      RECT 1.52 0.395 1.96 0.725 ;
  END
END scs130lp_o2bb2a_0

MACRO scs130lp_o2bb2a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2a_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.21 1.38 2.165 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.55 1.755 2 2.14 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 1.92 3.685 2.21 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.01 1.11 3.755 1.75 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 0.255 0.355 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.935 -0.085 3.265 0.545 ;
        RECT 0.525 -0.085 0.875 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.325 2.51 3.655 3.415 ;
        RECT 1.97 2.65 2.3 3.415 ;
        RECT 0.525 2.505 1.265 3.415 ;
        RECT 0.525 1.815 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.54 0.715 3.695 0.885 ;
      RECT 3.435 0.28 3.695 0.885 ;
      RECT 2.54 0.28 2.765 0.885 ;
      RECT 2.505 2.65 2.84 2.92 ;
      RECT 2.67 1.055 2.84 2.92 ;
      RECT 0.525 0.86 0.865 1.515 ;
      RECT 2.175 1.055 2.84 1.225 ;
      RECT 2.175 0.28 2.37 1.225 ;
      RECT 0.525 0.86 1.32 1.03 ;
      RECT 1.045 0.28 1.32 1.03 ;
      RECT 2.075 0.28 2.37 0.62 ;
      RECT 1.045 0.28 2.37 0.53 ;
      RECT 1.435 2.35 1.675 2.835 ;
      RECT 2.24 1.405 2.5 2.48 ;
      RECT 1.485 2.31 2.5 2.48 ;
      RECT 1.55 1.405 2.5 1.575 ;
      RECT 1.55 0.7 1.88 1.575 ;
  END
END scs130lp_o2bb2a_1

MACRO scs130lp_o2bb2a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2a_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 0.47 3.235 1.515 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 0.345 2.3 1.095 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.42 0.995 0.84 1.665 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 0.995 1.295 1.665 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.915 0.255 4.185 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.355 -0.085 4.605 1.095 ;
        RECT 3.405 -0.085 3.745 1.015 ;
        RECT 0.745 -0.085 1.075 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.355 1.815 4.605 3.415 ;
        RECT 3.375 2.025 3.745 3.415 ;
        RECT 1.825 2.095 2.155 3.415 ;
        RECT 0.295 1.835 0.625 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.325 2.665 3.205 2.835 ;
      RECT 3.035 1.685 3.205 2.835 ;
      RECT 2.325 1.755 2.495 2.835 ;
      RECT 1.14 1.835 1.655 2.515 ;
      RECT 1.465 1.755 2.495 1.925 ;
      RECT 3.035 1.685 3.745 1.855 ;
      RECT 3.495 1.185 3.745 1.855 ;
      RECT 1.465 0.995 1.645 2.515 ;
      RECT 1.465 0.995 1.895 1.165 ;
      RECT 1.66 0.28 1.895 1.165 ;
      RECT 2.665 0.28 2.855 2.485 ;
      RECT 1.815 1.335 2.855 1.585 ;
      RECT 2.47 0.28 2.855 1.585 ;
      RECT 0.295 0.655 1.49 0.825 ;
      RECT 1.245 0.28 1.49 0.825 ;
      RECT 0.295 0.28 0.575 0.825 ;
  END
END scs130lp_o2bb2a_2

MACRO scs130lp_o2bb2a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2a_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.92 1.085 5.17 1.515 ;
        RECT 3.645 1.085 5.17 1.255 ;
        RECT 3.645 1.085 4.175 1.515 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.345 1.425 4.75 1.76 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.845 1.345 2.095 1.65 ;
        RECT 0.625 2.31 2.025 2.5 ;
        RECT 1.845 1.345 2.025 2.5 ;
        RECT 0.625 1.405 0.815 2.5 ;
        RECT 0.33 1.405 0.815 1.645 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.405 1.315 1.76 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.68 1.745 7.595 1.925 ;
        RECT 7.345 1.045 7.595 1.925 ;
        RECT 5.875 1.045 7.595 1.235 ;
        RECT 6.805 0.255 6.995 1.235 ;
        RECT 6.54 1.745 6.72 3.075 ;
        RECT 5.875 0.255 6.135 1.235 ;
        RECT 5.68 1.745 5.87 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 7.165 -0.085 7.495 0.875 ;
        RECT 6.305 -0.085 6.635 0.875 ;
        RECT 5.175 -0.085 5.705 0.915 ;
        RECT 3.385 -0.085 3.645 0.555 ;
        RECT 1.495 -0.085 1.825 0.485 ;
        RECT 0.635 -0.085 0.965 0.895 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.9 2.095 7.23 3.415 ;
        RECT 6.04 2.095 6.37 3.415 ;
        RECT 5.105 2.78 5.435 3.415 ;
        RECT 4.23 2.78 4.56 3.415 ;
        RECT 3.03 2.78 3.7 3.415 ;
        RECT 1.935 2.67 2.42 3.415 ;
        RECT 2.195 1.795 2.42 3.415 ;
        RECT 0.205 1.815 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.59 1.73 2.86 3.075 ;
      RECT 2.59 2.43 5.51 2.61 ;
      RECT 5.34 1.405 5.51 2.61 ;
      RECT 2.59 1.73 2.93 2.61 ;
      RECT 0.985 1.93 1.665 2.14 ;
      RECT 1.485 0.995 1.665 2.14 ;
      RECT 2.59 0.605 2.76 3.075 ;
      RECT 5.34 1.405 7.175 1.575 ;
      RECT 1.485 0.995 2.76 1.175 ;
      RECT 2.505 0.605 2.76 1.175 ;
      RECT 4.745 0.255 5.005 0.915 ;
      RECT 3.815 0.255 5.005 0.485 ;
      RECT 3.295 1.93 4.945 2.26 ;
      RECT 3.295 0.725 3.475 2.26 ;
      RECT 2.93 1.185 3.475 1.515 ;
      RECT 3.295 0.725 4.575 0.915 ;
      RECT 4.245 0.655 4.575 0.915 ;
      RECT 0.205 1.065 1.315 1.235 ;
      RECT 1.135 0.255 1.315 1.235 ;
      RECT 0.205 0.255 0.465 1.235 ;
      RECT 2.93 0.255 3.125 1.015 ;
      RECT 1.135 0.655 2.335 0.825 ;
      RECT 2.005 0.255 2.335 0.825 ;
      RECT 1.135 0.255 1.325 0.825 ;
      RECT 2.005 0.255 3.125 0.435 ;
      RECT 0.625 2.67 1.765 3 ;
  END
END scs130lp_o2bb2a_4

MACRO scs130lp_o2bb2a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2a_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.55 1.315 2.15 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.21 2.275 1.88 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.65 1.55 4.22 1.88 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.55 3.41 1.88 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.265 0.455 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.445 -0.085 3.695 1.02 ;
        RECT 0.915 -0.085 1.245 0.68 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.875 2.06 4.205 3.415 ;
        RECT 2.025 2.84 2.355 3.415 ;
        RECT 0.655 2.84 0.985 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.015 1.2 4.205 1.37 ;
      RECT 3.875 0.85 4.205 1.37 ;
      RECT 3.015 0.69 3.265 1.37 ;
      RECT 2.815 2.06 3.145 3.065 ;
      RECT 0.635 2.49 3.145 2.66 ;
      RECT 0.635 0.86 0.805 2.66 ;
      RECT 0.635 0.86 0.965 1.19 ;
      RECT 2.505 0.775 2.835 1.15 ;
      RECT 0.635 0.86 2.835 1.03 ;
      RECT 1.735 0.265 2.065 0.68 ;
      RECT 1.735 0.265 2.835 0.595 ;
      RECT 1.495 2.06 2.625 2.31 ;
      RECT 2.455 1.5 2.625 2.31 ;
      RECT 2.455 1.5 2.785 1.83 ;
  END
END scs130lp_o2bb2a_lp

MACRO scs130lp_o2bb2a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2a_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.925 1.115 2.49 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.47 1.655 1.38 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.265 1.58 3.685 2.515 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.58 2.975 2.49 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.345 0.5 0.675 ;
        RECT 0.155 2.655 0.39 2.985 ;
        RECT 0.155 0.345 0.325 2.985 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.86 -0.085 3.19 1.045 ;
        RECT 0.72 -0.085 0.93 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.13 2.845 3.46 3.415 ;
        RECT 1.695 2.845 2.025 3.415 ;
        RECT 0.57 2.845 0.9 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.47 1.225 3.58 1.395 ;
      RECT 3.37 0.945 3.58 1.395 ;
      RECT 2.47 0.945 2.68 1.395 ;
      RECT 2.205 2.67 2.61 3 ;
      RECT 2.205 1.575 2.375 3 ;
      RECT 0.505 1.575 2.375 1.745 ;
      RECT 2.04 0.945 2.25 1.745 ;
      RECT 0.505 0.935 0.675 1.745 ;
      RECT 1.08 2.67 1.515 3 ;
      RECT 1.345 2.265 1.515 3 ;
      RECT 1.345 2.265 2.025 2.435 ;
      RECT 1.695 1.925 2.025 2.435 ;
      RECT 1.835 0.275 2.425 0.605 ;
  END
END scs130lp_o2bb2a_m

MACRO scs130lp_o2bb2ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2ai_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.825 0.39 2.96 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 0.825 1.005 2.195 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.89 1.12 3.275 2.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.12 2.49 1.825 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2905 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 2.005 2.305 3.065 ;
        RECT 1.555 2.005 2.305 2.175 ;
        RECT 1.555 1.57 1.895 2.175 ;
        RECT 1.725 0.28 1.895 2.175 ;
        RECT 1.545 0.28 1.895 0.61 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.475 -0.085 2.735 0.61 ;
        RECT 0.13 -0.085 0.46 0.655 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.795 2.395 3.125 3.415 ;
        RECT 1.555 2.395 1.865 3.415 ;
        RECT 0.685 2.395 0.98 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.065 0.78 3.205 0.95 ;
      RECT 2.905 0.28 3.205 0.95 ;
      RECT 2.065 0.28 2.305 0.95 ;
      RECT 1.15 2.395 1.385 3.065 ;
      RECT 1.195 0.81 1.385 3.065 ;
      RECT 1.195 0.81 1.545 1.4 ;
      RECT 1.195 0.325 1.365 3.065 ;
      RECT 0.95 0.325 1.365 0.655 ;
  END
END scs130lp_o2bb2ai_0

MACRO scs130lp_o2bb2ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2ai_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.45 1.75 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.21 1.035 1.54 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.185 3.275 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.185 2.735 2.995 ;
        RECT 2.33 1.185 2.735 1.585 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6762 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.99 1.755 2.335 3.075 ;
        RECT 1.93 1.065 2.1 1.925 ;
        RECT 1.545 1.065 2.1 1.235 ;
        RECT 1.545 0.255 1.785 1.235 ;
        RECT 1.525 0.255 1.785 0.65 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.455 -0.085 2.785 0.555 ;
        RECT 0.12 -0.085 0.45 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.915 1.92 3.245 3.415 ;
        RECT 0.98 2.095 1.82 3.415 ;
        RECT 0.12 1.92 0.45 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.27 0.725 3.245 1.015 ;
      RECT 2.975 0.265 3.245 1.015 ;
      RECT 1.955 0.285 2.285 0.895 ;
      RECT 0.62 1.755 0.81 3.075 ;
      RECT 0.62 1.755 1.415 1.925 ;
      RECT 1.205 1.405 1.415 1.925 ;
      RECT 1.205 1.405 1.76 1.675 ;
      RECT 1.205 0.82 1.375 1.925 ;
      RECT 0.985 0.255 1.315 1.04 ;
  END
END scs130lp_o2bb2ai_1

MACRO scs130lp_o2bb2ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2ai_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.92 2.01 2.09 ;
        RECT 1.695 1.295 2.01 2.09 ;
        RECT 0.085 1.375 0.805 2.09 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.21 1.455 1.75 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.565 1.92 5.675 2.09 ;
        RECT 5.325 1.295 5.675 2.09 ;
        RECT 3.565 1.345 3.815 2.09 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.995 1.21 5.155 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9912 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.9 2.26 4.55 2.59 ;
        RECT 2.9 0.595 3.23 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 4.7 -0.085 5.03 0.7 ;
        RECT 3.84 -0.085 4.17 0.7 ;
        RECT 1.89 -0.085 2.22 0.66 ;
        RECT 0.17 -0.085 0.475 1.205 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 5.13 2.26 5.46 3.415 ;
        RECT 3.4 2.76 3.63 3.415 ;
        RECT 1.925 2.62 2.73 3.415 ;
        RECT 2.52 1.815 2.73 3.415 ;
        RECT 1.03 2.6 1.36 3.415 ;
        RECT 0.17 2.27 0.5 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.52 0.255 2.73 1.205 ;
      RECT 3.41 0.87 5.46 1.04 ;
      RECT 5.2 0.325 5.46 1.04 ;
      RECT 4.34 0.325 4.53 1.04 ;
      RECT 3.41 0.255 3.67 1.04 ;
      RECT 2.52 0.255 3.67 0.425 ;
      RECT 3.8 2.76 4.95 3.075 ;
      RECT 4.72 2.26 4.95 3.075 ;
      RECT 1.53 2.26 1.755 3.075 ;
      RECT 0.67 2.26 0.86 3.075 ;
      RECT 1.53 2.26 2.35 2.45 ;
      RECT 2.18 0.83 2.35 2.45 ;
      RECT 0.67 2.26 2.35 2.43 ;
      RECT 2.18 1.375 2.565 1.625 ;
      RECT 1.03 0.83 2.35 1.04 ;
      RECT 0.645 0.305 0.86 1.09 ;
      RECT 0.645 0.305 1.71 0.66 ;
  END
END scs130lp_o2bb2ai_2

MACRO scs130lp_o2bb2ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2ai_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.905 1.425 7.935 1.595 ;
        RECT 5.905 1.21 6.565 1.595 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.285 1.425 9.635 1.595 ;
        RECT 8.285 1.17 8.975 1.595 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.055 1.95 3.81 2.13 ;
        RECT 3.48 1.425 3.81 2.13 ;
        RECT 1.055 1.425 1.415 2.13 ;
        RECT 0.405 1.425 1.415 1.645 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.425 3.205 1.78 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9656 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.995 1.075 5.515 1.245 ;
        RECT 5.185 0.615 5.515 1.245 ;
        RECT 5.075 1.775 5.265 3.075 ;
        RECT 3.995 1.775 5.265 1.945 ;
        RECT 4.165 0.605 4.495 1.245 ;
        RECT 4.215 1.775 4.405 3.075 ;
        RECT 2.015 2.3 4.405 2.63 ;
        RECT 3.995 1.775 4.405 2.63 ;
        RECT 3.995 1.075 4.165 2.63 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 7.425 -0.085 7.755 0.905 ;
        RECT 6.565 -0.085 6.895 0.7 ;
        RECT 3.145 -0.085 3.485 0.915 ;
        RECT 2.285 -0.085 2.615 0.905 ;
        RECT 1.425 -0.085 1.755 0.905 ;
        RECT 0.565 -0.085 0.895 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.56 2.115 9.89 3.415 ;
        RECT 8.7 2.125 9.03 3.415 ;
        RECT 7.5 2.125 8.17 3.415 ;
        RECT 6.64 2.125 6.97 3.415 ;
        RECT 5.435 2.125 6.11 3.415 ;
        RECT 4.575 2.115 4.905 3.415 ;
        RECT 3.745 2.8 4.045 3.415 ;
        RECT 1.065 2.69 1.395 3.415 ;
        RECT 0.265 1.815 0.475 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.21 1.765 9.39 3.075 ;
      RECT 8.34 1.765 8.53 3.075 ;
      RECT 7.14 1.765 7.33 3.075 ;
      RECT 6.28 1.765 6.47 3.075 ;
      RECT 5.555 1.765 9.995 1.945 ;
      RECT 9.815 1.075 9.995 1.945 ;
      RECT 5.555 1.425 5.725 1.945 ;
      RECT 4.345 1.425 5.725 1.595 ;
      RECT 9.145 1.075 9.995 1.255 ;
      RECT 9.145 0.605 9.475 1.255 ;
      RECT 8.285 0.815 9.475 1 ;
      RECT 8.285 0.605 8.585 1 ;
      RECT 7.055 1.075 8.115 1.245 ;
      RECT 7.925 0.265 8.115 1.245 ;
      RECT 7.055 0.87 7.255 1.245 ;
      RECT 7.065 0.305 7.255 1.245 ;
      RECT 6.135 0.87 7.255 1.04 ;
      RECT 9.655 0.265 9.985 0.905 ;
      RECT 6.135 0.305 6.395 1.04 ;
      RECT 8.755 0.265 8.975 0.635 ;
      RECT 7.925 0.265 9.985 0.435 ;
      RECT 0.135 1.085 3.825 1.255 ;
      RECT 3.655 0.265 3.825 1.255 ;
      RECT 0.135 1.075 2.975 1.255 ;
      RECT 2.785 0.305 2.975 1.255 ;
      RECT 1.925 0.305 2.115 1.255 ;
      RECT 1.065 0.305 1.255 1.255 ;
      RECT 0.135 0.305 0.385 1.255 ;
      RECT 5.685 0.265 5.945 1.04 ;
      RECT 3.655 0.265 3.985 0.905 ;
      RECT 4.675 0.265 5.005 0.895 ;
      RECT 3.655 0.265 5.945 0.435 ;
      RECT 1.575 2.8 3.575 3.075 ;
      RECT 0.695 2.35 0.895 3.075 ;
      RECT 1.575 2.35 1.785 3.075 ;
      RECT 0.695 2.35 1.785 2.52 ;
      RECT 0.695 1.815 0.885 3.075 ;
  END
END scs130lp_o2bb2ai_4

MACRO scs130lp_o2bb2ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2ai_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.49 1.895 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.02 0.905 1.315 1.575 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.895 1.185 3.26 1.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.265 1.185 2.725 1.78 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3997 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.895 2.115 2.225 3.065 ;
        RECT 1.925 1.255 2.095 3.065 ;
        RECT 1.545 1.255 2.095 1.425 ;
        RECT 1.545 0.395 1.875 1.425 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.405 -0.085 2.735 0.675 ;
        RECT 0.115 -0.085 0.445 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.915 2.075 3.245 3.415 ;
        RECT 1.23 2.115 1.56 3.415 ;
        RECT 0.16 2.075 0.49 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.055 0.845 3.195 1.015 ;
      RECT 2.915 0.46 3.195 1.015 ;
      RECT 2.055 0.46 2.225 1.015 ;
      RECT 0.67 1.765 1.03 3.065 ;
      RECT 0.67 1.765 1.755 1.935 ;
      RECT 1.505 1.605 1.755 1.935 ;
      RECT 0.67 0.555 0.84 3.065 ;
      RECT 0.67 0.555 1.265 0.725 ;
      RECT 0.935 0.265 1.265 0.725 ;
  END
END scs130lp_o2bb2ai_lp

MACRO scs130lp_o2bb2ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o2bb2ai_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.955 0.355 2.49 ;
        RECT 0.155 0.84 0.325 2.49 ;
    END
  END A1N
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 1.04 2.12 ;
    END
  END A2N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.84 1.21 3.205 2.49 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.245 2.12 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2289 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.655 2.32 2.245 2.49 ;
        RECT 1.655 0.5 1.865 2.49 ;
        RECT 1.495 2.715 1.825 2.925 ;
        RECT 1.655 0.5 1.825 2.925 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.515 -0.085 2.725 0.68 ;
        RECT 0.125 -0.085 0.455 0.655 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.285 2.845 2.615 3.415 ;
        RECT 0.975 2.845 1.305 3.415 ;
        RECT 0.095 2.845 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.085 0.86 3.155 1.03 ;
      RECT 2.945 0.5 3.155 1.03 ;
      RECT 2.085 0.52 2.295 1.03 ;
      RECT 0.605 2.345 0.795 2.985 ;
      RECT 0.605 2.345 1.44 2.515 ;
      RECT 1.27 0.45 1.44 2.515 ;
      RECT 0.915 0.45 1.44 0.66 ;
  END
END scs130lp_o2bb2ai_m

MACRO scs130lp_o311a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311a_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1 1.36 1.865 ;
        RECT 1.025 0.84 1.335 1.865 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.195 1.85 1.865 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.02 1.08 2.35 1.835 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.52 1.115 2.92 1.865 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.475 0.82 3.755 1.86 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4237 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.32 0.81 0.65 ;
        RECT 0.085 2.385 0.67 3.065 ;
        RECT 0.085 0.32 0.38 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.865 -0.085 2.195 0.57 ;
        RECT 0.985 -0.085 1.315 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.74 2.395 3.07 3.415 ;
        RECT 0.84 2.385 1.17 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.24 2.045 3.515 3.065 ;
      RECT 2.24 2.045 2.57 3.065 ;
      RECT 0.55 2.045 3.515 2.215 ;
      RECT 3.09 0.32 3.305 2.215 ;
      RECT 0.55 1.545 0.855 2.215 ;
      RECT 3.09 0.32 3.485 0.65 ;
      RECT 1.505 0.74 2.695 0.91 ;
      RECT 2.365 0.32 2.695 0.91 ;
      RECT 1.505 0.32 1.695 0.91 ;
  END
END scs130lp_o311a_0

MACRO scs130lp_o311a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311a_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.185 1.345 1.515 ;
        RECT 1.085 0.38 1.285 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 1.185 1.875 1.435 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.185 2.335 1.515 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.185 2.875 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.425 1.195 3.75 1.525 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.095 2.045 0.67 3.075 ;
        RECT 0.095 0.255 0.365 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.885 -0.085 2.215 0.675 ;
        RECT 0.585 -0.085 0.915 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.8 2.045 3.13 3.415 ;
        RECT 0.84 2.045 1.17 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.38 1.705 3.65 3.075 ;
      RECT 2.26 1.705 2.59 3.075 ;
      RECT 0.535 1.705 3.65 1.875 ;
      RECT 3.075 0.255 3.245 1.875 ;
      RECT 0.535 1.345 0.795 1.875 ;
      RECT 3.075 0.255 3.62 1.015 ;
      RECT 1.455 0.845 2.78 1.015 ;
      RECT 2.45 0.255 2.78 1.015 ;
      RECT 1.455 0.255 1.675 1.015 ;
  END
END scs130lp_o311a_1

MACRO scs130lp_o311a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311a_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.345 1.83 2.96 ;
        RECT 1.445 1.345 1.83 1.685 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 1.345 2.305 2.96 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 1.345 2.81 1.735 ;
        RECT 2.475 1.345 2.725 2.96 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.98 1.345 3.315 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.845 1.335 4.235 1.76 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.695 0.915 3.075 ;
        RECT 0.595 0.255 0.81 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 2.345 -0.085 2.675 0.495 ;
        RECT 0.98 -0.085 1.65 0.835 ;
        RECT 0.12 -0.085 0.425 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.305 2.27 3.635 3.415 ;
        RECT 1.155 1.855 1.425 3.415 ;
        RECT 0.155 1.815 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.805 1.93 4.065 3.075 ;
      RECT 2.895 1.92 3.135 3.075 ;
      RECT 2.895 1.93 4.065 2.1 ;
      RECT 2.895 1.92 3.675 2.1 ;
      RECT 3.485 1.005 3.675 2.1 ;
      RECT 0.98 1.005 1.235 1.515 ;
      RECT 0.98 1.005 3.675 1.175 ;
      RECT 3.52 0.255 4.06 1.165 ;
      RECT 1.82 0.665 3.215 0.835 ;
      RECT 2.885 0.255 3.215 0.835 ;
      RECT 1.82 0.255 2.15 0.835 ;
  END
END scs130lp_o311a_2

MACRO scs130lp_o311a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311a_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.285 1.425 8.075 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.85 1.425 7.115 1.76 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.955 1.21 5.68 1.515 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 1.195 3.785 1.525 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.965 1.195 3.265 1.525 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.835 1.755 2.025 3.075 ;
        RECT 0.085 1.755 2.025 1.925 ;
        RECT 0.085 1.065 1.69 1.235 ;
        RECT 1.46 0.255 1.69 1.235 ;
        RECT 0.975 1.755 1.165 3.075 ;
        RECT 0.085 1.055 0.79 1.235 ;
        RECT 0.6 0.255 0.79 1.235 ;
        RECT 0.085 1.055 0.36 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.23 -0.085 7.56 0.915 ;
        RECT 6.37 -0.085 6.7 0.915 ;
        RECT 5.01 -0.085 5.84 0.7 ;
        RECT 1.86 -0.085 2.15 1.105 ;
        RECT 0.96 -0.085 1.29 0.895 ;
        RECT 0.1 -0.085 0.43 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.23 2.27 7.56 3.415 ;
        RECT 3.99 2.045 4.32 3.415 ;
        RECT 3.095 2.045 3.425 3.415 ;
        RECT 2.195 2.045 2.525 3.415 ;
        RECT 1.335 2.105 1.665 3.415 ;
        RECT 0.475 2.095 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6 1.085 7.99 1.255 ;
      RECT 7.73 0.255 7.99 1.255 ;
      RECT 6.87 0.255 7.06 1.255 ;
      RECT 6 0.87 6.2 1.255 ;
      RECT 6.01 0.255 6.2 1.255 ;
      RECT 3.955 0.87 6.2 1.04 ;
      RECT 3.63 0.615 3.96 1.025 ;
      RECT 3.63 0.855 4.84 1.025 ;
      RECT 4.58 0.255 4.84 1.04 ;
      RECT 7.73 1.93 7.99 3.075 ;
      RECT 6.87 1.93 7.06 3.075 ;
      RECT 5.94 1.93 6.2 2.735 ;
      RECT 5.94 1.93 7.99 2.1 ;
      RECT 4.51 2.905 6.7 3.075 ;
      RECT 6.37 2.27 6.7 3.075 ;
      RECT 5.405 1.705 5.68 3.075 ;
      RECT 4.51 2.045 4.84 3.075 ;
      RECT 3.595 1.705 3.82 3.075 ;
      RECT 2.695 1.705 2.925 3.075 ;
      RECT 5.01 1.705 5.235 2.735 ;
      RECT 2.195 1.705 5.235 1.875 ;
      RECT 2.195 1.405 2.795 1.875 ;
      RECT 0.53 1.405 2.795 1.585 ;
      RECT 2.32 0.765 2.795 1.875 ;
      RECT 2.32 0.765 3.1 1.015 ;
      RECT 3.27 0.255 3.46 1.025 ;
      RECT 4.13 0.255 4.39 0.685 ;
      RECT 2.34 0.255 3.46 0.595 ;
      RECT 2.34 0.255 4.39 0.435 ;
  END
END scs130lp_o311a_4

MACRO scs130lp_o311a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311a_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.99 1.55 1.32 1.92 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.55 1.86 1.92 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.55 2.36 1.88 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.53 1.55 2.86 1.92 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.03 1.55 3.41 1.92 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 2.115 0.46 3.065 ;
        RECT 0.1 0.44 0.445 1.085 ;
        RECT 0.1 0.44 0.27 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.85 -0.085 2.18 1.02 ;
        RECT 0.905 -0.085 1.155 1.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.835 2.45 3.165 3.415 ;
        RECT 0.66 2.45 0.99 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.455 2.1 3.75 3.065 ;
      RECT 3.58 0.74 3.75 3.065 ;
      RECT 2.295 2.1 2.625 3.065 ;
      RECT 0.64 2.1 3.75 2.27 ;
      RECT 0.64 1.265 0.81 2.27 ;
      RECT 0.45 1.265 0.81 1.935 ;
      RECT 3.15 0.74 3.75 1.07 ;
      RECT 1.5 1.2 2.69 1.37 ;
      RECT 2.36 0.685 2.69 1.37 ;
      RECT 1.5 0.685 1.67 1.37 ;
      RECT 1.34 0.685 1.67 1.145 ;
  END
END scs130lp_o311a_lp

MACRO scs130lp_o311a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311a_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 1.105 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 1.155 1.765 2.49 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.96 1.075 2.29 1.585 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.795 2.75 1.465 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 0.84 3.685 2.49 ;
    END
  END C1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.231 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.33 0.635 0.66 ;
        RECT 0.155 1.965 0.41 2.295 ;
        RECT 0.155 0.33 0.325 2.295 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.715 -0.085 1.925 0.545 ;
        RECT 0.855 -0.085 1.065 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.685 2.115 2.895 3.415 ;
        RECT 0.59 2.155 0.92 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.025 2.855 2.355 3.025 ;
      RECT 2.145 1.765 2.355 3.025 ;
      RECT 3.115 1.765 3.305 2.275 ;
      RECT 3.135 0.405 3.305 2.275 ;
      RECT 2.145 1.765 3.305 1.935 ;
      RECT 3.135 0.405 3.495 0.615 ;
      RECT 1.285 0.725 2.335 0.895 ;
      RECT 2.145 0.345 2.335 0.895 ;
      RECT 1.285 0.345 1.495 0.895 ;
  END
END scs130lp_o311a_m

MACRO scs130lp_o311ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311ai_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.535 0.77 0.84 1.835 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 1.16 1.355 1.83 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.16 1.865 1.78 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.16 2.495 1.78 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 0.84 3.275 1.78 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4985 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.705 1.95 3.275 2.99 ;
        RECT 2.665 0.285 3.01 0.615 ;
        RECT 2.665 0.285 2.835 2.12 ;
        RECT 1.705 1.95 3.275 2.12 ;
        RECT 1.705 1.95 2.035 2.98 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.43 -0.085 1.715 0.615 ;
        RECT 0.51 -0.085 0.84 0.6 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.205 2.32 2.535 3.415 ;
        RECT 0.51 2.32 0.84 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.01 0.785 2.19 0.99 ;
      RECT 1.885 0.285 2.19 0.99 ;
      RECT 1.01 0.285 1.26 0.99 ;
  END
END scs130lp_o311ai_0

MACRO scs130lp_o311ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311ai_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.345 0.86 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 1.345 1.355 2.98 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.345 1.865 1.775 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.345 2.405 1.78 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 1.21 3.275 1.77 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0479 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.91 1.94 3.275 3.075 ;
        RECT 2.575 0.255 3.24 1.04 ;
        RECT 1.795 1.95 3.275 2.12 ;
        RECT 2.575 1.94 3.275 2.12 ;
        RECT 2.575 0.255 2.765 2.12 ;
        RECT 1.795 1.95 2.125 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.31 -0.085 1.64 0.835 ;
        RECT 0.41 -0.085 0.67 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.38 2.29 2.71 3.415 ;
        RECT 0.41 1.92 0.74 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.84 1.005 2.405 1.175 ;
      RECT 1.81 0.265 2.405 1.175 ;
      RECT 0.84 0.265 1.14 1.175 ;
  END
END scs130lp_o311ai_1

MACRO scs130lp_o311ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311ai_2 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.185 0.945 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.185 1.9 1.435 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.34 1.185 3.205 1.525 ;
        RECT 2.07 1.185 3.205 1.435 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.47 1.185 4.285 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.295 1.21 5.675 1.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8186 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.405 1.715 5.665 3.075 ;
        RECT 4.455 0.87 5.665 1.04 ;
        RECT 5.395 0.335 5.665 1.04 ;
        RECT 4.545 1.715 5.665 1.885 ;
        RECT 2.375 1.695 5.125 1.865 ;
        RECT 4.545 0.87 5.125 1.885 ;
        RECT 4.455 0.595 4.805 1.865 ;
        RECT 4.545 0.595 4.735 3.075 ;
        RECT 3.305 1.695 3.495 3.075 ;
        RECT 2.375 1.695 2.635 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.76 0.085 ;
        RECT 2.325 -0.085 3 0.675 ;
        RECT 1.425 -0.085 1.755 0.675 ;
        RECT 0.565 -0.085 0.895 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.76 3.415 ;
        RECT 4.905 2.055 5.235 3.415 ;
        RECT 3.665 2.035 4.375 3.415 ;
        RECT 0.565 1.945 0.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.975 0.255 5.225 0.7 ;
      RECT 3.525 0.255 3.855 0.675 ;
      RECT 3.525 0.255 5.225 0.425 ;
      RECT 0.135 0.845 4.285 1.015 ;
      RECT 4.025 0.595 4.285 1.015 ;
      RECT 3.17 0.255 3.355 1.015 ;
      RECT 1.925 0.255 2.155 1.015 ;
      RECT 1.065 0.255 1.255 1.015 ;
      RECT 0.135 0.255 0.395 1.015 ;
      RECT 1.425 2.905 3.135 3.075 ;
      RECT 2.805 2.035 3.135 3.075 ;
      RECT 1.425 1.945 1.755 3.075 ;
      RECT 1.065 1.605 1.255 3.075 ;
      RECT 0.135 1.605 0.395 3.075 ;
      RECT 1.925 1.605 2.185 2.735 ;
      RECT 0.135 1.605 2.185 1.775 ;
  END
END scs130lp_o311ai_2

MACRO scs130lp_o311ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311ai_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.09 1.18 1.86 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 1.18 3.795 1.435 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.465 1.425 6.095 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.265 1.425 7.615 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.785 1.425 9.995 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.0618 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.31 1.92 9.57 3.075 ;
        RECT 4.08 1.085 9.43 1.255 ;
        RECT 9.1 0.595 9.43 1.255 ;
        RECT 4.08 1.92 9.57 2.09 ;
        RECT 8.45 1.92 8.64 3.075 ;
        RECT 8.1 0.595 8.43 1.255 ;
        RECT 7.59 1.92 7.78 3.075 ;
        RECT 6.73 1.92 6.92 3.075 ;
        RECT 4.08 1.92 6.92 2.12 ;
        RECT 5.87 1.92 6.06 3.075 ;
        RECT 5.01 1.92 5.2 2.735 ;
        RECT 4.08 1.92 4.34 2.735 ;
        RECT 4.08 1.085 4.295 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 5.27 -0.085 5.6 0.555 ;
        RECT 4.41 -0.085 4.74 0.575 ;
        RECT 3.55 -0.085 3.88 0.575 ;
        RECT 2.69 -0.085 3.02 0.67 ;
        RECT 1.83 -0.085 2.16 0.67 ;
        RECT 0.97 -0.085 1.3 0.67 ;
        RECT 0.11 -0.085 0.44 1.01 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.81 2.26 9.14 3.415 ;
        RECT 7.95 2.26 8.28 3.415 ;
        RECT 7.09 2.26 7.42 3.415 ;
        RECT 6.23 2.29 6.56 3.415 ;
        RECT 1.4 1.945 1.73 3.415 ;
        RECT 0.54 1.945 0.87 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.6 0.255 9.86 1.19 ;
      RECT 8.6 0.255 8.93 0.915 ;
      RECT 7.6 0.255 7.93 0.915 ;
      RECT 5.81 0.255 7.93 0.555 ;
      RECT 5.81 0.255 9.86 0.425 ;
      RECT 0.61 0.84 3.91 1.01 ;
      RECT 4.91 0.725 7.43 0.915 ;
      RECT 3.19 0.745 7.43 0.915 ;
      RECT 2.33 0.255 2.52 1.01 ;
      RECT 1.47 0.255 1.66 1.01 ;
      RECT 0.61 0.255 0.8 1.01 ;
      RECT 4.05 0.255 4.24 0.915 ;
      RECT 3.19 0.255 3.38 1.01 ;
      RECT 4.91 0.255 5.1 0.915 ;
      RECT 2.26 2.905 5.7 3.075 ;
      RECT 5.37 2.29 5.7 3.075 ;
      RECT 4.51 2.29 4.84 3.075 ;
      RECT 3.12 1.945 3.45 3.075 ;
      RECT 2.26 1.945 2.59 3.075 ;
      RECT 1.9 1.605 2.09 3.075 ;
      RECT 1.04 1.605 1.23 3.075 ;
      RECT 0.11 1.605 0.37 3.075 ;
      RECT 3.62 1.605 3.88 2.735 ;
      RECT 2.76 1.605 2.95 2.735 ;
      RECT 0.11 1.605 3.88 1.775 ;
  END
END scs130lp_o311ai_4

MACRO scs130lp_o311ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311ai_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.115 1.295 0.445 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.88 1.605 1.315 2.89 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.3 2.275 0.67 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.605 2.275 2.15 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.47 1.365 2.8 1.78 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6847 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.725 2.075 3.235 3.065 ;
        RECT 3.005 0.44 3.235 3.065 ;
        RECT 2.595 0.72 3.235 1.18 ;
        RECT 1.645 2.33 3.235 2.5 ;
        RECT 1.645 2.33 1.975 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.055 -0.085 1.385 1.075 ;
        RECT 0.115 -0.085 0.445 1.115 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.175 2.68 2.505 3.415 ;
        RECT 0.115 2.075 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.625 1.255 2.055 1.425 ;
      RECT 1.725 0.85 2.055 1.425 ;
      RECT 0.625 0.72 0.875 1.425 ;
  END
END scs130lp_o311ai_lp

MACRO scs130lp_o311ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o311ai_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.455 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 2.69 0.935 3.025 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 2.69 1.765 3.025 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.58 2.245 1.75 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.955 2.725 1.75 ;
        RECT 2.555 0.84 2.725 1.75 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3402 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 1.93 2.725 2.325 ;
        RECT 2.175 0.45 2.635 0.66 ;
        RECT 1.495 1.93 2.725 2.1 ;
        RECT 0.635 1.21 2.345 1.38 ;
        RECT 2.175 0.45 2.345 1.38 ;
        RECT 0.635 2.32 1.705 2.49 ;
        RECT 1.495 1.93 1.705 2.49 ;
        RECT 0.635 1.21 0.805 2.49 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.085 -0.085 1.415 0.66 ;
        RECT 0.225 -0.085 0.555 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.945 2.28 2.275 3.415 ;
        RECT 0.235 2.125 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.735 0.84 1.785 1.01 ;
      RECT 1.595 0.52 1.785 1.01 ;
      RECT 0.735 0.52 0.905 1.01 ;
  END
END scs130lp_o311ai_m

MACRO scs130lp_o31a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31a_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.08 1.35 1.865 ;
        RECT 1.015 0.82 1.295 1.865 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.08 1.81 1.865 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.98 1.195 2.35 1.865 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.52 1.055 2.92 1.865 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.32 0.595 0.65 ;
        RECT 0.085 2.385 0.57 3.075 ;
        RECT 0.085 0.32 0.35 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.855 -0.085 2.185 0.545 ;
        RECT 0.825 -0.085 1.155 0.65 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.615 2.385 2.945 3.415 ;
        RECT 0.815 2.385 1.145 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.115 2.035 2.445 3.055 ;
      RECT 0.53 2.035 3.275 2.215 ;
      RECT 3.09 0.32 3.275 2.215 ;
      RECT 0.53 1.545 0.845 2.215 ;
      RECT 2.775 0.32 3.275 0.65 ;
      RECT 1.465 0.715 2.605 0.885 ;
      RECT 2.355 0.32 2.605 0.885 ;
      RECT 1.465 0.32 1.685 0.885 ;
      RECT 1.365 0.32 1.685 0.65 ;
  END
END scs130lp_o31a_0

MACRO scs130lp_o31a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31a_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.21 1.285 1.755 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 1.345 1.835 1.76 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.345 2.375 1.76 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.345 2.925 1.76 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.255 0.385 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.87 -0.085 2.2 0.835 ;
        RECT 0.555 -0.085 1.25 1.025 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.79 2.27 3.12 3.415 ;
        RECT 0.555 2.27 1.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.29 1.93 2.62 3.075 ;
      RECT 0.555 1.93 3.275 2.1 ;
      RECT 3.095 0.255 3.275 2.1 ;
      RECT 0.555 1.195 0.805 2.1 ;
      RECT 2.825 0.255 3.275 1.105 ;
      RECT 1.455 1.005 2.655 1.175 ;
      RECT 2.37 0.255 2.655 1.175 ;
      RECT 1.455 0.255 1.7 1.175 ;
  END
END scs130lp_o31a_1

MACRO scs130lp_o31a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31a_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.375 1.815 2.945 ;
        RECT 1.445 1.375 1.815 1.675 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.985 1.375 2.315 2.945 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.345 2.785 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.305 1.345 3.755 1.75 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 1.695 0.915 3.075 ;
        RECT 0.595 0.255 0.815 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.26 -0.085 2.59 0.495 ;
        RECT 0.985 -0.085 1.59 0.865 ;
        RECT 0.12 -0.085 0.395 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.295 1.92 3.515 3.415 ;
        RECT 1.105 1.82 1.355 3.415 ;
        RECT 0.155 1.815 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.71 1.93 3.125 3.075 ;
      RECT 2.955 1.005 3.125 3.075 ;
      RECT 0.985 1.035 1.235 1.515 ;
      RECT 0.985 1.035 1.93 1.205 ;
      RECT 3.26 0.255 3.52 1.175 ;
      RECT 1.76 1.005 3.52 1.175 ;
      RECT 1.76 0.665 3.09 0.835 ;
      RECT 2.76 0.255 3.09 0.835 ;
      RECT 1.76 0.255 2.09 0.835 ;
  END
END scs130lp_o31a_2

MACRO scs130lp_o31a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31a_4 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.375 1.21 6.095 1.535 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.92 1.705 6.595 1.875 ;
        RECT 6.265 1.295 6.595 1.875 ;
        RECT 4.85 1.345 5.205 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.515 1.425 4.68 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.425 3.335 2.12 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.795 1.755 1.975 3.075 ;
        RECT 0.085 1.755 1.975 1.925 ;
        RECT 0.085 1.055 1.75 1.225 ;
        RECT 1.56 0.255 1.75 1.225 ;
        RECT 0.925 1.755 1.115 3.075 ;
        RECT 0.7 0.255 0.89 1.225 ;
        RECT 0.085 1.055 0.335 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.72 0.085 ;
        RECT 5.865 -0.085 6.195 0.7 ;
        RECT 4.925 -0.085 5.255 0.7 ;
        RECT 3.99 -0.085 4.32 0.895 ;
        RECT 1.92 -0.085 2.25 1.105 ;
        RECT 1.06 -0.085 1.39 0.885 ;
        RECT 0.2 -0.085 0.53 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.72 3.415 ;
        RECT 6.365 2.435 6.625 3.415 ;
        RECT 5.425 2.435 6.625 2.665 ;
        RECT 3.005 2.63 3.335 3.415 ;
        RECT 2.145 1.815 2.475 3.415 ;
        RECT 1.285 2.095 1.615 3.415 ;
        RECT 0.425 2.095 0.755 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.63 1.075 4.71 1.245 ;
      RECT 4.49 0.305 4.71 1.245 ;
      RECT 3.63 0.255 3.82 1.245 ;
      RECT 4.49 0.87 6.625 1.04 ;
      RECT 6.365 0.305 6.625 1.04 ;
      RECT 2.62 0.255 2.95 0.905 ;
      RECT 5.435 0.305 5.695 1.04 ;
      RECT 4.49 0.305 4.75 1.04 ;
      RECT 2.62 0.255 3.82 0.435 ;
      RECT 4.43 1.92 4.75 3.075 ;
      RECT 4.43 2.045 6.625 2.265 ;
      RECT 3.56 1.92 4.75 2.12 ;
      RECT 4.925 2.835 6.195 3.075 ;
      RECT 4.925 2.435 5.255 3.075 ;
      RECT 3.99 2.29 4.26 3.075 ;
      RECT 2.645 1.075 2.825 3.075 ;
      RECT 2.645 2.29 4.26 2.46 ;
      RECT 2.645 1.075 2.835 2.46 ;
      RECT 0.505 1.405 2.835 1.575 ;
      RECT 2.635 1.075 2.835 1.575 ;
      RECT 2.635 1.075 3.46 1.245 ;
      RECT 3.13 0.605 3.46 1.245 ;
  END
END scs130lp_o31a_4

MACRO scs130lp_o31a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31a_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.17 2.39 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.17 1.85 1.84 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.125 1.315 1.795 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.125 0.805 1.795 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.925 1.92 3.27 3.065 ;
        RECT 3.1 0.265 3.27 3.065 ;
        RECT 2.915 0.265 3.27 0.725 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.125 -0.085 2.455 0.725 ;
        RECT 1.185 -0.085 1.515 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.315 2.37 2.645 3.415 ;
        RECT 0.195 2.325 0.525 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.725 1.975 1.055 3.065 ;
      RECT 0.725 2.02 2.745 2.19 ;
      RECT 2.575 0.93 2.745 2.19 ;
      RECT 0.09 1.975 1.055 2.145 ;
      RECT 0.09 0.265 0.26 2.145 ;
      RECT 2.575 0.93 2.92 1.6 ;
      RECT 0.09 0.265 0.495 0.725 ;
      RECT 0.675 0.775 1.945 0.945 ;
      RECT 1.695 0.265 1.945 0.945 ;
      RECT 0.675 0.265 1.005 0.945 ;
  END
END scs130lp_o31a_lp

MACRO scs130lp_o31a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31a_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.945 1.155 1.285 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.485 1.155 1.765 2.49 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 1.015 2.275 1.525 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.47 2.735 1.435 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.675 0.58 2.235 ;
        RECT 0.37 0.345 0.58 2.235 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.62 -0.085 1.95 0.485 ;
        RECT 0.8 -0.085 1.01 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.61 2.155 2.94 3.415 ;
        RECT 0.76 2.095 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.15 2.67 1.48 3.025 ;
      RECT 1.15 2.67 2.34 2.84 ;
      RECT 2.13 1.805 2.34 2.84 ;
      RECT 2.13 1.805 3.105 1.975 ;
      RECT 2.915 0.345 3.105 1.975 ;
      RECT 1.23 0.665 2.375 0.835 ;
      RECT 2.185 0.345 2.375 0.835 ;
      RECT 1.23 0.345 1.44 0.835 ;
  END
END scs130lp_o31a_m

MACRO scs130lp_o31ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31ai_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.41 2.225 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.58 1.13 1.005 2.225 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.36 1.105 1.895 1.81 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 0.84 2.255 1.81 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4333 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.485 1.98 2.79 2.225 ;
        RECT 2.425 0.34 2.79 2.225 ;
        RECT 2.065 0.34 2.79 0.67 ;
        RECT 1.485 1.98 1.815 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.145 -0.085 1.475 0.595 ;
        RECT 0.235 -0.085 0.565 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.985 2.395 2.245 3.415 ;
        RECT 0.275 2.395 0.605 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.735 0.765 1.895 0.935 ;
      RECT 1.645 0.37 1.895 0.935 ;
      RECT 0.735 0.37 0.975 0.935 ;
  END
END scs130lp_o31ai_0

MACRO scs130lp_o31ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31ai_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.395 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.565 1.345 1.01 1.75 ;
        RECT 0.595 1.345 0.87 2.99 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.375 2.255 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.425 1.375 2.795 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0227 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.18 1.035 2.555 1.205 ;
        RECT 2.295 0.255 2.555 1.205 ;
        RECT 1.04 1.95 2.11 3.075 ;
        RECT 1.18 1.035 1.35 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 0.945 -0.085 1.625 0.525 ;
        RECT 0.095 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.28 1.92 2.54 3.415 ;
        RECT 0.095 1.92 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.595 0.695 0.855 1.095 ;
      RECT 0.595 0.695 2.125 0.865 ;
      RECT 1.795 0.265 2.125 0.865 ;
      RECT 0.595 0.255 0.775 1.095 ;
  END
END scs130lp_o31ai_1

MACRO scs130lp_o31ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31ai_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 1.285 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.455 1.21 2.275 1.525 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 1.425 3.415 1.755 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.645 1.415 4.715 1.585 ;
        RECT 4.26 1.21 4.715 1.585 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4511 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 1.755 4.705 3.075 ;
        RECT 3.595 1.755 4.705 1.925 ;
        RECT 2.685 1.075 4.08 1.245 ;
        RECT 3.75 0.595 4.08 1.245 ;
        RECT 3.415 1.925 3.775 3.075 ;
        RECT 2.42 1.925 3.775 2.12 ;
        RECT 2.685 1.075 2.855 2.12 ;
        RECT 2.42 1.815 2.75 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 2.82 -0.085 3.15 0.565 ;
        RECT 1.58 -0.085 2.175 0.7 ;
        RECT 0.68 -0.085 1.01 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.945 2.095 4.275 3.415 ;
        RECT 0.68 2.035 0.87 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.25 0.255 4.51 1.04 ;
      RECT 0.25 0.87 2.515 1.04 ;
      RECT 3.32 0.255 3.58 0.905 ;
      RECT 2.345 0.735 3.58 0.905 ;
      RECT 1.18 0.315 1.41 1.04 ;
      RECT 0.25 0.315 0.51 1.04 ;
      RECT 2.345 0.285 2.65 0.905 ;
      RECT 3.32 0.255 4.51 0.425 ;
      RECT 1.54 2.905 3.18 3.075 ;
      RECT 2.92 2.29 3.18 3.075 ;
      RECT 1.54 2.035 1.73 3.075 ;
      RECT 1.04 1.695 1.37 3.075 ;
      RECT 0.18 1.695 0.51 3.075 ;
      RECT 1.9 1.695 2.23 2.735 ;
      RECT 0.18 1.695 2.23 1.865 ;
  END
END scs130lp_o31ai_2

MACRO scs130lp_o31ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31ai_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.94 1.425 2.29 1.595 ;
        RECT 1.485 1.425 1.835 1.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.46 1.325 3.67 1.505 ;
        RECT 2.46 1.075 2.985 1.505 ;
        RECT 0.33 1.075 2.985 1.245 ;
        RECT 0.33 1.075 0.66 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.11 1.335 7.72 1.535 ;
        RECT 3.985 1.695 7.28 1.865 ;
        RECT 7.11 1.335 7.28 1.865 ;
        RECT 3.985 1.325 5.005 1.865 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.24 1.345 6.93 1.525 ;
        RECT 5.435 1.2 6.575 1.525 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.3184 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.46 1.705 8.075 1.875 ;
        RECT 7.89 0.995 8.075 1.875 ;
        RECT 6.745 0.995 8.075 1.165 ;
        RECT 7.335 2.035 7.63 2.715 ;
        RECT 7.46 1.705 7.63 2.715 ;
        RECT 5.005 2.035 7.63 2.24 ;
        RECT 5.465 0.7 6.925 1.03 ;
        RECT 5.005 2.035 5.185 2.725 ;
        RECT 4.145 2.035 7.63 2.215 ;
        RECT 4.145 2.035 4.335 2.735 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.605 -0.085 7.935 0.825 ;
        RECT 4.55 -0.085 4.88 0.805 ;
        RECT 3.645 -0.085 3.975 0.805 ;
        RECT 2.785 -0.085 3.115 0.565 ;
        RECT 1.925 -0.085 2.255 0.565 ;
        RECT 1.065 -0.085 1.395 0.565 ;
        RECT 0.205 -0.085 0.465 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 6.555 2.75 6.825 3.415 ;
        RECT 5.695 2.75 5.905 3.415 ;
        RECT 1.995 2.61 2.185 3.415 ;
        RECT 1.135 2.61 1.325 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.645 2.905 5.525 3.075 ;
      RECT 5.355 2.41 5.525 3.075 ;
      RECT 0.205 1.815 0.465 3.075 ;
      RECT 6.995 2.895 8.06 3.065 ;
      RECT 7.8 2.045 8.06 3.065 ;
      RECT 4.505 2.895 5.525 3.075 ;
      RECT 3.645 2.035 3.975 3.075 ;
      RECT 6.995 2.41 7.165 3.065 ;
      RECT 4.505 2.385 4.835 3.075 ;
      RECT 2.855 1.815 3.075 2.715 ;
      RECT 5.355 2.41 7.165 2.58 ;
      RECT 1.145 1.93 2.175 2.1 ;
      RECT 3.645 1.705 3.815 3.075 ;
      RECT 2.005 1.815 3.075 1.985 ;
      RECT 0.205 1.815 1.315 1.985 ;
      RECT 2.865 1.705 3.815 1.875 ;
      RECT 3.275 0.985 5.265 1.155 ;
      RECT 5.065 0.255 5.265 1.155 ;
      RECT 4.155 0.425 4.38 1.155 ;
      RECT 3.275 0.735 3.475 1.155 ;
      RECT 3.285 0.255 3.475 1.155 ;
      RECT 0.635 0.735 3.475 0.905 ;
      RECT 7.095 0.255 7.425 0.825 ;
      RECT 2.425 0.255 2.615 0.905 ;
      RECT 1.565 0.255 1.755 0.905 ;
      RECT 0.635 0.255 0.895 0.905 ;
      RECT 5.065 0.255 7.425 0.53 ;
      RECT 2.355 2.885 3.475 3.075 ;
      RECT 3.245 2.055 3.475 3.075 ;
      RECT 1.495 2.27 1.825 3.075 ;
      RECT 0.635 2.155 0.965 3.075 ;
      RECT 2.355 2.155 2.685 3.075 ;
      RECT 0.635 2.27 2.685 2.44 ;
  END
END scs130lp_o31ai_4

MACRO scs130lp_o31ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31ai_lp 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.11 0.55 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.925 1.265 1.315 2.89 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.225 1.825 1.895 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.225 2.395 1.895 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4733 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 2.29 2.755 2.52 ;
        RECT 2.585 0.265 2.755 2.52 ;
        RECT 2.31 0.265 2.755 0.725 ;
        RECT 1.565 2.075 2.05 3.065 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.29 -0.085 1.62 0.695 ;
        RECT 0.27 -0.085 0.6 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 2.29 2.7 2.62 3.415 ;
        RECT 0.13 2.075 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.78 0.875 2.13 1.045 ;
      RECT 1.8 0.265 2.13 1.045 ;
      RECT 0.78 0.265 1.11 1.045 ;
  END
END scs130lp_o31ai_lp

MACRO scs130lp_o31ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o31ai_m 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.175 0.47 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.88 1.535 1.285 2.49 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.535 1.765 2.205 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.285 2.245 0.64 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2625 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 2.435 2.305 2.605 ;
        RECT 1.975 0.835 2.305 2.605 ;
        RECT 1.525 2.69 1.765 3.02 ;
        RECT 1.595 2.435 1.765 3.02 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.095 -0.085 1.285 0.935 ;
        RECT 0.235 -0.085 0.445 0.955 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.955 2.785 2.165 3.415 ;
        RECT 0.315 2.845 0.645 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.665 1.115 1.795 1.285 ;
      RECT 1.465 0.835 1.795 1.285 ;
      RECT 0.665 0.775 0.875 1.285 ;
  END
END scs130lp_o31ai_m

MACRO scs130lp_o32a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32a_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.84 1.285 1.855 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.48 1.185 1.845 1.855 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 1.185 2.355 1.855 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.425 0.955 3.755 2.12 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.185 2.895 1.855 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.395 0.69 3.065 ;
        RECT 0.085 0.47 0.6 0.8 ;
        RECT 0.085 0.47 0.385 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.87 -0.085 2.2 0.675 ;
        RECT 0.83 -0.085 1.16 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.16 2.395 3.49 3.415 ;
        RECT 0.92 2.385 1.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.465 0.845 2.68 1.015 ;
      RECT 2.41 0.255 2.68 1.015 ;
      RECT 1.465 0.385 1.66 1.015 ;
      RECT 3.415 0.255 3.67 0.785 ;
      RECT 1.33 0.385 1.66 0.67 ;
      RECT 2.41 0.255 3.67 0.425 ;
      RECT 2.31 2.025 2.64 3.075 ;
      RECT 0.555 2.025 3.255 2.215 ;
      RECT 3.065 0.845 3.255 2.215 ;
      RECT 0.555 1.545 0.815 2.215 ;
      RECT 2.91 0.595 3.245 0.855 ;
  END
END scs130lp_o32a_0

MACRO scs130lp_o32a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32a_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.07 1.21 1.355 1.755 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.21 1.845 1.76 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 1.21 2.37 1.76 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.44 1.21 3.755 2.12 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.54 1.345 2.92 1.76 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.325 0.6 1.175 ;
        RECT 0.085 1.815 0.56 3.075 ;
        RECT 0.085 0.325 0.265 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.655 -0.085 2.325 0.7 ;
        RECT 0.77 -0.085 1.1 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.355 2.29 3.685 3.415 ;
        RECT 0.8 2.27 1.13 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.43 0.255 3.71 1.04 ;
      RECT 1.27 0.87 2.73 1.04 ;
      RECT 2.495 0.255 2.73 1.04 ;
      RECT 1.27 0.305 1.485 1.04 ;
      RECT 2.495 0.255 3.71 0.425 ;
      RECT 2.215 1.93 2.91 3.075 ;
      RECT 0.73 1.93 3.26 2.1 ;
      RECT 3.09 0.595 3.26 2.1 ;
      RECT 0.73 1.345 0.9 2.1 ;
      RECT 0.44 1.345 0.9 1.645 ;
      RECT 2.9 0.595 3.26 1.175 ;
  END
END scs130lp_o32a_1

MACRO scs130lp_o32a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32a_2 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.185 1.815 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.985 1.21 2.315 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.485 1.21 2.855 1.515 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.845 1.21 4.235 1.83 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 1.21 3.315 1.54 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.585 0.255 0.81 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 2.25 -0.085 2.58 0.7 ;
        RECT 1.11 -0.085 1.44 1.035 ;
        RECT 0.12 -0.085 0.415 1.09 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.81 2 4.06 3.415 ;
        RECT 0.98 2.025 1.65 3.415 ;
        RECT 0.12 1.815 0.415 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.825 0.255 4.095 1.04 ;
      RECT 1.91 0.87 3.13 1.04 ;
      RECT 2.83 0.255 3.13 1.04 ;
      RECT 1.68 0.255 2.01 1.015 ;
      RECT 2.83 0.255 4.095 0.425 ;
      RECT 2.7 1.71 3.03 3.075 ;
      RECT 2.7 1.71 3.655 1.925 ;
      RECT 3.485 0.595 3.655 1.925 ;
      RECT 1.175 1.685 2.915 1.855 ;
      RECT 1.175 1.34 1.345 1.855 ;
      RECT 0.985 1.34 1.345 1.67 ;
      RECT 3.3 0.595 3.655 0.935 ;
  END
END scs130lp_o32a_2

MACRO scs130lp_o32a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32a_4 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 1.21 1.83 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.01 1.27 2.375 1.535 ;
        RECT 0.085 1.695 2.18 1.865 ;
        RECT 2.01 1.27 2.18 1.865 ;
        RECT 0.085 1.425 1.33 1.865 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 3.69 1.535 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 1.21 4.775 1.525 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.86 1.695 5.625 1.865 ;
        RECT 4.945 1.425 5.625 1.865 ;
        RECT 3.86 1.355 4.195 1.865 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.485 1.755 8.075 1.925 ;
        RECT 7.81 1.055 8.075 1.925 ;
        RECT 6.485 1.055 8.075 1.225 ;
        RECT 7.345 1.755 7.535 3.075 ;
        RECT 7.345 0.255 7.525 1.225 ;
        RECT 6.485 1.755 6.675 3.075 ;
        RECT 6.485 0.255 6.665 1.225 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.705 -0.085 8.035 0.885 ;
        RECT 6.845 -0.085 7.175 0.885 ;
        RECT 5.985 -0.085 6.315 0.905 ;
        RECT 2.73 -0.085 3.06 0.7 ;
        RECT 1.81 -0.085 2.14 0.7 ;
        RECT 0.61 -0.085 1.235 0.7 ;
        RECT 0.61 -0.085 0.94 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.705 2.095 8.035 3.415 ;
        RECT 6.845 2.095 7.175 3.415 ;
        RECT 5.985 2.375 6.315 3.415 ;
        RECT 4.525 2.715 4.855 3.415 ;
        RECT 1.38 2.715 1.71 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.455 2.035 5.715 3.075 ;
      RECT 2.71 2.905 3.92 3.075 ;
      RECT 3.66 2.035 3.92 3.075 ;
      RECT 2.71 2.045 3.04 3.075 ;
      RECT 3.66 2.035 6.3 2.205 ;
      RECT 5.795 1.075 6.3 2.205 ;
      RECT 5.795 1.395 7.64 1.585 ;
      RECT 4.955 1.075 6.3 1.255 ;
      RECT 4.025 0.595 4.275 1.185 ;
      RECT 4.955 0.615 5.285 1.255 ;
      RECT 4.025 0.87 5.285 1.04 ;
      RECT 4.025 0.595 4.355 1.04 ;
      RECT 0.18 1.085 1.33 1.255 ;
      RECT 1.16 0.87 1.33 1.255 ;
      RECT 0.18 0.305 0.44 1.255 ;
      RECT 1.16 0.87 3.855 1.04 ;
      RECT 3.23 0.255 3.855 1.04 ;
      RECT 5.465 0.255 5.795 0.895 ;
      RECT 2.31 0.305 2.56 1.04 ;
      RECT 1.405 0.255 1.64 1.04 ;
      RECT 4.525 0.255 4.785 0.7 ;
      RECT 4.525 0.255 5.795 0.435 ;
      RECT 3.23 0.255 5.795 0.425 ;
      RECT 5.025 2.375 5.285 3.075 ;
      RECT 4.09 2.375 4.355 3.075 ;
      RECT 4.09 2.375 5.285 2.545 ;
      RECT 2.35 1.705 2.54 3.075 ;
      RECT 0.52 2.035 0.78 3.065 ;
      RECT 3.21 1.705 3.47 2.735 ;
      RECT 0.52 2.035 2.54 2.205 ;
      RECT 2.35 1.705 3.47 1.875 ;
      RECT 1.88 2.375 2.18 3.075 ;
      RECT 0.95 2.375 1.21 3.075 ;
      RECT 0.95 2.375 2.18 2.545 ;
  END
END scs130lp_o32a_4

MACRO scs130lp_o32a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32a_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.515 1.395 2.845 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.975 1.33 2.305 1.78 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.435 1.395 1.795 1.78 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.18 0.435 1.78 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.615 1.425 1.225 2.89 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.375 1.92 3.735 3.065 ;
        RECT 3.565 0.425 3.735 3.065 ;
        RECT 3.395 0.425 3.735 0.885 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.605 -0.085 2.935 0.8 ;
        RECT 1.665 -0.085 1.995 0.45 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.835 2.31 3.165 3.415 ;
        RECT 0.185 2.075 0.435 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.405 1.96 1.655 3.065 ;
      RECT 1.405 1.96 3.195 2.13 ;
      RECT 3.025 0.98 3.195 2.13 ;
      RECT 3.025 1.07 3.385 1.74 ;
      RECT 0.645 0.98 3.195 1.15 ;
      RECT 0.645 0.615 0.975 1.15 ;
      RECT 0.135 0.265 0.465 0.945 ;
      RECT 1.155 0.63 2.425 0.8 ;
      RECT 2.175 0.425 2.425 0.8 ;
      RECT 1.155 0.265 1.485 0.8 ;
      RECT 0.135 0.265 1.485 0.435 ;
  END
END scs130lp_o32a_lp

MACRO scs130lp_o32a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32a_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.84 1.12 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.535 1.185 1.765 2.49 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.185 2.245 2.49 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.395 0.84 3.685 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.535 1.185 2.865 1.695 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.125 0.395 2.86 ;
        RECT 0.155 0.47 0.395 0.8 ;
        RECT 0.155 0.47 0.325 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 1.67 -0.085 2 0.655 ;
        RECT 0.575 -0.085 0.905 0.655 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.2 2.225 3.53 3.415 ;
        RECT 0.575 2.185 0.905 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.3 0.835 2.55 1.005 ;
      RECT 2.36 0.265 2.55 1.005 ;
      RECT 1.3 0.515 1.49 1.005 ;
      RECT 3.24 0.265 3.57 0.655 ;
      RECT 2.36 0.265 3.57 0.435 ;
      RECT 2.11 2.855 2.635 3.025 ;
      RECT 2.465 1.875 2.635 3.025 ;
      RECT 2.425 2.125 2.635 3.025 ;
      RECT 2.465 1.875 3.215 2.045 ;
      RECT 3.045 0.835 3.215 2.045 ;
      RECT 2.73 0.615 3.06 1.005 ;
  END
END scs130lp_o32a_m

MACRO scs130lp_o32ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32ai_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.21 2.955 2.22 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.21 2.335 2.95 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.555 1.21 1.835 2.95 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.455 2.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.56 1.355 2.23 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4158 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 2.435 1.385 3.075 ;
        RECT 0.625 2.435 1.385 2.95 ;
        RECT 0.625 0.595 0.955 1.39 ;
        RECT 0.625 0.595 0.815 2.95 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.8 -0.085 3.07 0.785 ;
        RECT 1.485 -0.085 2.21 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.62 2.445 2.83 3.415 ;
        RECT 0.205 2.435 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.125 0.87 2.58 1.04 ;
      RECT 2.38 0.455 2.58 1.04 ;
      RECT 1.125 0.255 1.315 1.04 ;
      RECT 0.125 0.255 0.455 0.67 ;
      RECT 0.125 0.255 1.315 0.425 ;
  END
END scs130lp_o32ai_0

MACRO scs130lp_o32ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32ai_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.21 3.275 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.21 2.725 1.83 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.21 1.865 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.935 0.605 1.75 ;
        RECT 0.085 0.84 0.6 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.345 1.415 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1466 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.775 1.92 1.87 3.075 ;
        RECT 0.775 0.595 1.1 1.175 ;
        RECT 0.775 0.595 0.945 3.075 ;
        RECT 0.77 0.595 1.1 0.765 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.9 -0.085 3.23 1.04 ;
        RECT 1.7 -0.085 2.37 0.7 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.87 1.92 3.2 3.415 ;
        RECT 0.34 1.92 0.605 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.27 0.87 2.73 1.04 ;
      RECT 2.54 0.325 2.73 1.04 ;
      RECT 1.27 0.255 1.53 1.04 ;
      RECT 0.34 0.255 0.6 0.67 ;
      RECT 0.34 0.255 1.53 0.425 ;
  END
END scs130lp_o32ai_1

MACRO scs130lp_o32ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32ai_2 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.815 1.21 6.155 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.505 1.21 4.645 1.525 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 1.415 2.835 1.75 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.425 1.83 1.75 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.425 1.295 1.75 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2432 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.075 3.335 2.735 ;
        RECT 0.585 1.92 3.335 2.09 ;
        RECT 0.585 1.075 3.335 1.245 ;
        RECT 1.605 0.595 1.935 1.245 ;
        RECT 0.585 1.92 0.915 2.735 ;
        RECT 0.585 0.595 0.915 1.245 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 4.835 -0.085 5.165 0.7 ;
        RECT 3.945 -0.085 4.275 0.7 ;
        RECT 2.615 -0.085 3.405 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.71 1.815 6.005 3.415 ;
        RECT 4.815 2.045 5.145 3.415 ;
        RECT 1.445 2.62 1.775 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.155 0.255 0.415 1.185 ;
      RECT 3.505 0.87 5.595 1.04 ;
      RECT 5.335 0.315 5.595 1.04 ;
      RECT 2.115 0.735 3.775 0.905 ;
      RECT 1.095 0.255 1.425 0.905 ;
      RECT 4.465 0.315 4.665 1.04 ;
      RECT 3.575 0.315 3.775 1.04 ;
      RECT 2.115 0.255 2.445 0.905 ;
      RECT 0.155 0.255 2.445 0.425 ;
      RECT 5.315 1.705 5.54 3.075 ;
      RECT 3.865 1.705 4.195 2.735 ;
      RECT 3.865 1.705 5.54 1.875 ;
      RECT 2.555 2.905 4.625 3.075 ;
      RECT 4.365 2.045 4.625 3.075 ;
      RECT 3.505 1.815 3.695 3.075 ;
      RECT 2.555 2.26 2.825 3.075 ;
      RECT 1.945 2.26 2.205 3.075 ;
      RECT 0.155 2.905 1.275 3.075 ;
      RECT 1.085 2.26 1.275 3.075 ;
      RECT 0.155 1.92 0.415 3.075 ;
      RECT 1.085 2.26 2.205 2.45 ;
  END
END scs130lp_o32ai_2

MACRO scs130lp_o32ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32ai_4 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.425 1.21 10.455 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.185 1.21 8.215 1.495 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.965 1.335 5.655 1.76 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.425 3.755 1.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.375 1.855 1.76 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.352 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.54 1.93 6.005 2.1 ;
        RECT 5.835 0.995 6.005 2.1 ;
        RECT 3.19 0.995 6.005 1.165 ;
        RECT 5.415 1.93 5.68 2.735 ;
        RECT 4.57 1.93 4.82 2.735 ;
        RECT 0.57 1.005 3.41 1.175 ;
        RECT 3.19 0.615 3.38 1.175 ;
        RECT 2.33 0.595 2.52 1.175 ;
        RECT 1.4 1.93 1.765 2.735 ;
        RECT 1.47 0.595 1.66 1.175 ;
        RECT 0.54 1.93 0.87 2.735 ;
        RECT 0.57 0.595 0.8 1.175 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.41 -0.085 9.74 0.7 ;
        RECT 8.55 -0.085 8.88 0.7 ;
        RECT 7.31 -0.085 7.94 0.7 ;
        RECT 6.405 -0.085 6.745 0.475 ;
        RECT 5.09 -0.085 5.42 0.485 ;
        RECT 4.09 -0.085 4.42 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.88 1.815 10.17 3.415 ;
        RECT 8.98 2.005 9.31 3.415 ;
        RECT 8.12 2.005 8.45 3.415 ;
        RECT 3.155 2.62 3.485 3.415 ;
        RECT 2.295 2.62 2.625 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.11 0.255 0.4 1.095 ;
      RECT 6.175 0.87 10.17 1.04 ;
      RECT 9.91 0.255 10.17 1.04 ;
      RECT 9.05 0.255 9.24 1.04 ;
      RECT 8.11 0.255 8.38 1.04 ;
      RECT 6.915 0.255 7.14 1.04 ;
      RECT 6.175 0.645 6.345 1.04 ;
      RECT 2.69 0.255 3.02 0.835 ;
      RECT 1.83 0.255 2.16 0.835 ;
      RECT 0.97 0.255 1.3 0.835 ;
      RECT 3.55 0.655 6.345 0.825 ;
      RECT 5.59 0.255 6.235 0.825 ;
      RECT 4.59 0.255 4.92 0.825 ;
      RECT 3.55 0.255 3.88 0.825 ;
      RECT 2.69 0.255 3.88 0.445 ;
      RECT 0.11 0.255 3.88 0.425 ;
      RECT 9.48 1.665 9.71 3.075 ;
      RECT 8.62 1.665 8.81 3.075 ;
      RECT 7.145 1.665 7.41 2.735 ;
      RECT 6.29 1.665 6.545 2.735 ;
      RECT 6.29 1.665 9.71 1.835 ;
      RECT 4.105 2.905 7.875 3.075 ;
      RECT 7.58 2.005 7.875 3.075 ;
      RECT 6.715 2.005 6.975 3.075 ;
      RECT 5.85 2.27 6.12 3.075 ;
      RECT 4.99 2.27 5.245 3.075 ;
      RECT 4.105 2.27 4.375 3.075 ;
      RECT 3.655 2.27 3.915 3.075 ;
      RECT 2.795 2.27 2.985 3.075 ;
      RECT 0.11 2.905 2.125 3.075 ;
      RECT 1.935 2.27 2.125 3.075 ;
      RECT 1.04 2.27 1.23 3.075 ;
      RECT 0.11 1.94 0.37 3.075 ;
      RECT 1.935 2.27 3.915 2.45 ;
  END
END scs130lp_o32ai_4

MACRO scs130lp_o32ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32ai_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.915 1.295 3.245 1.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.605 2.395 2.89 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.605 1.825 2.89 ;
        RECT 1.495 1.605 1.825 1.935 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.515 0.605 1.845 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.265 1.795 1.04 ;
        RECT 0.93 0.265 1.795 0.555 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3976 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 2.115 1.385 3.065 ;
        RECT 1.085 1.92 1.315 3.065 ;
        RECT 0.785 1.92 1.315 2.09 ;
        RECT 0.785 1.085 0.955 2.09 ;
        RECT 0.625 1.085 0.955 1.335 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.915 -0.085 3.245 1.115 ;
        RECT 1.975 -0.085 2.225 1.075 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.86 2.075 3.19 3.415 ;
        RECT 0.115 2.075 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.135 1.255 2.735 1.425 ;
      RECT 2.405 0.745 2.735 1.425 ;
      RECT 0.115 0.735 0.445 1.335 ;
      RECT 1.135 0.735 1.385 1.425 ;
      RECT 0.115 0.735 1.385 0.905 ;
  END
END scs130lp_o32ai_lp

MACRO scs130lp_o32ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o32ai_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.89 0.84 3.205 2.49 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.21 2.255 2.49 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.21 1.765 2.49 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.49 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 1.21 1.285 2.49 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2352 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 2.67 2.725 3 ;
        RECT 0.8 0.62 1.13 1.01 ;
        RECT 0.655 0.84 0.825 3 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.56 -0.085 2.89 0.66 ;
        RECT 1.68 -0.085 2.01 0.64 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.905 2.785 3.095 3.415 ;
        RECT 0.265 2.785 0.455 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.31 0.82 2.38 0.99 ;
      RECT 2.19 0.52 2.38 0.99 ;
      RECT 1.31 0.27 1.5 0.99 ;
      RECT 0.29 0.27 0.62 0.66 ;
      RECT 0.29 0.27 1.5 0.44 ;
  END
END scs130lp_o32ai_m

MACRO scs130lp_o41a_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41a_0 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.405 1.035 3.735 2.18 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.945 1.14 3.205 2.86 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.465 1.14 2.775 2.86 ;
        RECT 2.405 1.14 2.775 2.205 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.14 2.235 2.21 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.08 1.345 1.85 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 2.395 0.54 3.065 ;
        RECT 0.085 0.265 0.355 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.9 -0.085 3.23 0.525 ;
        RECT 2.035 -0.085 2.315 0.63 ;
        RECT 0.525 -0.085 0.855 0.57 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.375 2.395 3.69 3.415 ;
        RECT 0.71 2.395 1.04 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.61 0.8 2.7 0.97 ;
      RECT 3.4 0.3 3.705 0.865 ;
      RECT 2.485 0.695 3.705 0.865 ;
      RECT 1.61 0.3 1.865 0.97 ;
      RECT 2.485 0.3 2.73 0.865 ;
      RECT 1.21 2.395 1.99 3.075 ;
      RECT 1.21 2.045 1.425 3.075 ;
      RECT 0.525 2.045 1.425 2.215 ;
      RECT 0.525 0.74 0.775 2.215 ;
      RECT 0.525 0.74 1.44 0.91 ;
      RECT 1.14 0.3 1.44 0.91 ;
  END
END scs130lp_o41a_0

MACRO scs130lp_o41a_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41a_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.865 1.375 4.235 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.275 1.425 3.695 2.98 ;
        RECT 3.165 1.425 3.695 1.675 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.345 2.955 2.98 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.345 2.335 2.98 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.345 1.905 1.75 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2705 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.815 0.925 3.075 ;
        RECT 0.085 0.255 0.73 0.925 ;
        RECT 0.085 1.425 0.575 3.075 ;
        RECT 0.085 0.255 0.495 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.36 -0.085 3.69 0.835 ;
        RECT 2.35 -0.085 2.68 0.835 ;
        RECT 0.9 -0.085 1.23 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.865 1.92 4.16 3.415 ;
        RECT 1.155 2.27 1.485 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.88 1.005 4.16 1.175 ;
      RECT 3.86 0.255 4.16 1.175 ;
      RECT 2.86 0.255 3.19 1.175 ;
      RECT 1.88 0.255 2.15 1.175 ;
      RECT 1.655 1.925 1.905 3.075 ;
      RECT 1.255 1.925 1.905 2.1 ;
      RECT 1.255 0.995 1.425 2.1 ;
      RECT 0.78 1.095 1.425 1.525 ;
      RECT 0.9 0.995 1.425 1.525 ;
      RECT 1.42 0.255 1.71 1.165 ;
  END
END scs130lp_o41a_1

MACRO scs130lp_o41a_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41a_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.345 1.345 4.675 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.495 1.345 4.175 2.965 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.985 1.345 3.325 2.965 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.495 1.345 2.815 2.16 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.065 1.21 2.255 1.75 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 0.375 0.895 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.8 -0.085 4.13 0.835 ;
        RECT 2.83 -0.085 3.16 0.835 ;
        RECT 1.065 -0.085 1.395 1.175 ;
        RECT 0.205 -0.085 0.465 1.255 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 4.345 1.925 4.615 3.415 ;
        RECT 1.065 2.31 1.9 3.415 ;
        RECT 1.065 1.845 1.45 3.415 ;
        RECT 0.205 1.815 0.465 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.425 1.005 4.61 1.175 ;
      RECT 4.3 0.255 4.61 1.175 ;
      RECT 3.33 0.255 3.63 1.175 ;
      RECT 2.425 0.255 2.66 1.175 ;
      RECT 2.07 2.33 2.74 3.075 ;
      RECT 2.07 1.96 2.325 3.075 ;
      RECT 1.62 1.96 2.325 2.14 ;
      RECT 1.62 0.255 1.895 2.14 ;
      RECT 1.065 1.345 1.895 1.675 ;
      RECT 1.62 0.255 2.2 1.04 ;
  END
END scs130lp_o41a_2

MACRO scs130lp_o41a_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41a_4 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.395 1.21 7.595 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.345 1.21 6.225 1.435 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.985 1.21 5.175 1.435 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.455 1.21 3.815 1.435 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.69 1.21 3.285 1.435 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.47 1.755 1.66 3.075 ;
        RECT 0.085 1.055 1.66 1.225 ;
        RECT 1.47 0.255 1.66 1.225 ;
        RECT 0.085 1.755 1.66 1.925 ;
        RECT 0.61 1.755 0.8 3.075 ;
        RECT 0.61 0.255 0.8 1.225 ;
        RECT 0.085 1.055 0.335 1.925 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.755 -0.085 7.015 0.7 ;
        RECT 5.405 -0.085 6.15 0.7 ;
        RECT 4.545 -0.085 4.8 0.7 ;
        RECT 3.685 -0.085 3.945 0.7 ;
        RECT 1.83 -0.085 2.15 1.105 ;
        RECT 0.97 -0.085 1.3 0.885 ;
        RECT 0.11 -0.085 0.44 0.885 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.79 2.105 7.12 3.415 ;
        RECT 2.69 1.985 3.02 3.415 ;
        RECT 1.83 1.815 2.16 3.415 ;
        RECT 0.97 2.105 1.3 3.415 ;
        RECT 0.11 2.095 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.29 0.87 7.5 1.04 ;
      RECT 7.185 0.265 7.5 1.04 ;
      RECT 6.32 0.255 6.585 1.04 ;
      RECT 4.97 0.255 5.235 1.04 ;
      RECT 4.115 0.255 4.375 1.04 ;
      RECT 3.29 0.255 3.515 1.04 ;
      RECT 2.36 0.255 2.62 0.69 ;
      RECT 2.36 0.255 3.515 0.425 ;
      RECT 7.29 1.705 7.49 3.075 ;
      RECT 6.43 1.705 6.62 3.075 ;
      RECT 5.5 1.705 5.76 2.725 ;
      RECT 5.5 1.705 7.49 1.875 ;
      RECT 4.58 2.895 6.26 3.075 ;
      RECT 5.93 2.055 6.26 3.075 ;
      RECT 4.58 1.945 4.77 3.075 ;
      RECT 3.22 2.905 4.41 3.075 ;
      RECT 4.08 1.605 4.41 3.075 ;
      RECT 3.22 1.985 3.55 3.075 ;
      RECT 4.94 1.605 5.27 2.725 ;
      RECT 4.08 1.605 5.27 1.775 ;
      RECT 2.33 1.605 2.52 3.075 ;
      RECT 3.72 1.605 3.91 2.735 ;
      RECT 2.33 1.605 3.91 1.815 ;
      RECT 2.33 0.86 2.51 3.075 ;
      RECT 0.505 1.395 2.51 1.585 ;
      RECT 2.32 0.86 2.51 1.585 ;
      RECT 2.32 0.86 3.12 1.04 ;
      RECT 2.79 0.595 3.12 1.04 ;
  END
END scs130lp_o41a_4

MACRO scs130lp_o41a_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41a_lp 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.19 0.685 1.86 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.925 1.23 1.315 2.89 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.23 1.825 2.89 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.23 2.365 2.89 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.67 1.18 3.235 1.51 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.72 2.04 4.205 3.065 ;
        RECT 3.965 0.265 4.205 3.065 ;
        RECT 3.875 0.265 4.205 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.085 -0.085 3.415 0.65 ;
        RECT 1.665 -0.085 1.915 0.7 ;
        RECT 0.645 -0.085 0.975 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.075 2.04 3.405 3.415 ;
        RECT 0.13 2.04 0.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.545 1.69 2.875 3.065 ;
      RECT 2.545 1.69 3.745 1.86 ;
      RECT 3.415 1.19 3.745 1.86 ;
      RECT 3.415 0.83 3.585 1.86 ;
      RECT 2.525 0.83 3.585 1 ;
      RECT 2.525 0.265 2.855 1 ;
      RECT 1.155 0.88 2.345 1.05 ;
      RECT 2.095 0.265 2.345 1.05 ;
      RECT 0.135 0.84 1.485 1.01 ;
      RECT 1.155 0.265 1.485 1.05 ;
      RECT 0.135 0.265 0.465 1.01 ;
  END
END scs130lp_o41a_lp

MACRO scs130lp_o41a_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41a_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.37 1.21 3.685 2.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.21 2.89 2.49 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.145 2.32 2.49 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 1.765 2.86 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.955 1.21 1.285 2.265 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 2.795 0.62 3.005 ;
        RECT 0.155 0.345 0.365 3.005 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.825 -0.085 3.035 0.565 ;
        RECT 1.965 -0.085 2.175 0.565 ;
        RECT 0.585 -0.085 0.795 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.915 2.845 3.245 3.415 ;
        RECT 0.8 2.805 0.99 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.535 0.745 3.465 0.915 ;
      RECT 3.255 0.365 3.465 0.915 ;
      RECT 2.395 0.365 2.605 0.915 ;
      RECT 1.535 0.365 1.745 0.915 ;
      RECT 1.225 2.445 1.415 2.985 ;
      RECT 0.545 2.445 1.415 2.615 ;
      RECT 0.545 0.725 0.715 2.615 ;
      RECT 0.545 0.725 1.315 0.895 ;
      RECT 1.105 0.365 1.315 0.895 ;
  END
END scs130lp_o41a_m

MACRO scs130lp_o41ai_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41ai_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.915 1.17 3.275 2.19 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.27 1.17 2.745 2.235 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 2.045 2.06 3.025 ;
        RECT 1.595 1.17 2.06 3.025 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 1.205 1.425 1.875 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.595 0.815 0.895 1.85 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4879 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.03 2.055 1.33 3.065 ;
        RECT 0.1 2.055 1.33 2.225 ;
        RECT 0.1 0.315 0.93 0.645 ;
        RECT 0.1 0.315 0.415 2.225 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.48 -0.085 2.8 0.66 ;
        RECT 1.54 -0.085 1.87 0.66 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.71 2.405 3.085 3.415 ;
        RECT 0.57 2.405 0.86 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.1 0.83 3.265 1 ;
      RECT 2.97 0.33 3.265 1 ;
      RECT 2.04 0.33 2.31 1 ;
      RECT 1.1 0.33 1.37 1 ;
  END
END scs130lp_o41ai_0

MACRO scs130lp_o41ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41ai_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.21 3.275 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.03 1.425 2.4 2.965 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.53 1.425 1.86 2.965 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.07 1.345 1.36 1.78 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.375 0.455 1.75 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.865 1.95 1.165 3.075 ;
        RECT 0.73 1.345 0.9 2.17 ;
        RECT 0.625 1.025 0.795 1.515 ;
        RECT 0.085 0.255 0.635 1.195 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.255 -0.085 2.585 0.7 ;
        RECT 1.305 -0.085 1.635 0.835 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.695 1.925 3.065 3.415 ;
        RECT 0.31 2.34 0.695 3.415 ;
        RECT 0.31 1.925 0.56 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.965 1.005 2.735 1.175 ;
      RECT 2.755 0.255 3.085 1.04 ;
      RECT 1.805 0.87 3.085 1.04 ;
      RECT 0.965 0.255 1.135 1.175 ;
      RECT 1.805 0.255 2.085 1.175 ;
      RECT 0.805 0.255 1.135 0.855 ;
  END
END scs130lp_o41ai_1

MACRO scs130lp_o41ai_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41ai_2 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.32 1.335 6.115 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.93 1.335 5.15 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.385 1.335 3.76 1.75 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.455 1.335 3.215 1.75 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.015 1.065 1.525 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9408 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.955 1.335 2.285 2.715 ;
        RECT 0.615 1.705 2.285 1.875 ;
        RECT 1.235 1.335 2.285 1.875 ;
        RECT 1.235 0.595 1.485 1.875 ;
        RECT 0.615 1.705 0.835 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 4.83 -0.085 5.16 0.825 ;
        RECT 3.97 -0.085 4.3 0.825 ;
        RECT 3.07 -0.085 3.4 0.825 ;
        RECT 2.1 -0.085 2.43 0.825 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.29 2.26 5.62 3.415 ;
        RECT 1.005 2.045 1.335 3.415 ;
        RECT 0.145 1.815 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.79 1.92 6.05 3.075 ;
      RECT 4.93 1.92 5.12 3.075 ;
      RECT 4 1.92 4.26 2.735 ;
      RECT 4 1.92 6.05 2.09 ;
      RECT 1.655 0.995 5.61 1.165 ;
      RECT 5.34 0.255 5.61 1.165 ;
      RECT 4.47 0.255 4.66 1.165 ;
      RECT 3.57 0.255 3.8 1.165 ;
      RECT 2.62 0.255 2.9 1.165 ;
      RECT 1.655 0.255 1.925 1.165 ;
      RECT 0.735 0.255 1.065 0.845 ;
      RECT 0.735 0.255 1.925 0.425 ;
      RECT 3.05 2.905 4.76 3.075 ;
      RECT 4.43 2.26 4.76 3.075 ;
      RECT 3.05 2.26 3.38 3.075 ;
      RECT 1.525 2.895 2.84 3.075 ;
      RECT 2.51 1.92 2.84 3.075 ;
      RECT 1.525 2.045 1.785 3.075 ;
      RECT 3.55 1.92 3.81 2.735 ;
      RECT 2.51 1.92 3.81 2.09 ;
  END
END scs130lp_o41ai_2

MACRO scs130lp_o41ai_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41ai_4 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.765 1.21 10.475 1.525 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.745 1.345 8.435 1.525 ;
        RECT 6.745 1.345 7.335 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.845 1.345 6.575 1.75 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.985 1.355 4.255 1.525 ;
        RECT 2.985 1.355 3.685 1.76 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.375 2.815 1.76 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8816 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.02 1.705 4.675 1.875 ;
        RECT 4.425 1.015 4.675 1.875 ;
        RECT 1.385 1.015 4.675 1.185 ;
        RECT 4.02 1.705 4.35 2.725 ;
        RECT 0.99 1.93 4.35 2.1 ;
        RECT 3.16 1.93 3.49 2.725 ;
        RECT 2.28 0.595 2.47 1.185 ;
        RECT 1.86 1.93 2.04 3.075 ;
        RECT 1.385 0.595 1.61 1.185 ;
        RECT 0.99 1.93 1.18 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.66 -0.085 9.94 0.7 ;
        RECT 8.795 -0.085 9.07 0.7 ;
        RECT 7.84 -0.085 8.17 0.835 ;
        RECT 6.91 -0.085 7.24 0.835 ;
        RECT 6.05 -0.085 6.38 0.835 ;
        RECT 5.185 -0.085 5.515 0.835 ;
        RECT 4.17 -0.085 4.5 0.505 ;
        RECT 3.15 -0.085 3.48 0.505 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.7 2.045 10.03 3.415 ;
        RECT 8.84 2.045 9.17 3.415 ;
        RECT 2.21 2.27 2.54 3.415 ;
        RECT 1.35 2.27 1.68 3.415 ;
        RECT 0.49 1.93 0.82 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 10.2 1.695 10.46 3.075 ;
      RECT 9.34 1.695 9.53 3.075 ;
      RECT 8.48 1.695 8.67 3.075 ;
      RECT 6.69 1.92 6.95 2.685 ;
      RECT 7.62 1.695 7.88 2.49 ;
      RECT 6.69 1.92 7.88 2.1 ;
      RECT 7.62 1.695 10.46 1.875 ;
      RECT 4.845 1.005 8.585 1.175 ;
      RECT 0.92 0.255 1.215 1.095 ;
      RECT 10.11 0.255 10.39 1.04 ;
      RECT 8.34 0.87 10.39 1.04 ;
      RECT 7.41 0.255 7.67 1.175 ;
      RECT 6.55 0.255 6.74 1.175 ;
      RECT 5.69 0.255 5.88 1.175 ;
      RECT 4.845 0.255 5.015 1.175 ;
      RECT 9.24 0.255 9.49 1.04 ;
      RECT 8.34 0.255 8.625 1.04 ;
      RECT 2.64 0.675 5.015 0.845 ;
      RECT 4.68 0.255 5.015 0.845 ;
      RECT 1.78 0.255 2.11 0.845 ;
      RECT 3.66 0.255 3.99 0.845 ;
      RECT 2.64 0.255 2.97 0.845 ;
      RECT 0.92 0.255 2.97 0.425 ;
      RECT 4.88 2.855 8.31 3.075 ;
      RECT 8.05 2.045 8.31 3.075 ;
      RECT 7.12 2.735 8.31 3.075 ;
      RECT 5.74 2.395 6.07 3.075 ;
      RECT 4.88 2.395 5.21 3.075 ;
      RECT 7.12 2.27 7.45 3.075 ;
      RECT 2.73 2.895 4.71 3.075 ;
      RECT 4.52 2.045 4.71 3.075 ;
      RECT 3.66 2.27 3.85 3.075 ;
      RECT 2.73 2.27 2.99 3.075 ;
      RECT 6.24 1.92 6.5 2.685 ;
      RECT 5.38 1.92 5.57 2.685 ;
      RECT 4.52 2.045 6.5 2.225 ;
      RECT 4.845 1.92 6.5 2.225 ;
  END
END scs130lp_o41ai_4

MACRO scs130lp_o41ai_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41ai_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.81 1.225 3.235 1.895 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.055 1.265 2.445 2.89 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.545 1.265 1.875 2.89 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 1.125 1.335 1.795 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 1.125 0.825 1.795 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4333 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.74 1.975 1.07 3.065 ;
        RECT 0.115 1.975 1.07 2.145 ;
        RECT 0.115 0.265 0.56 0.725 ;
        RECT 0.115 0.265 0.285 2.145 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.32 -0.085 2.65 0.695 ;
        RECT 1.25 -0.085 1.58 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.91 2.075 3.24 3.415 ;
        RECT 0.21 2.325 0.54 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.81 0.875 3.16 1.045 ;
      RECT 2.83 0.265 3.16 1.045 ;
      RECT 0.74 0.775 2.14 0.945 ;
      RECT 1.81 0.265 2.14 1.045 ;
      RECT 0.74 0.265 1.07 0.945 ;
  END
END scs130lp_o41ai_lp

MACRO scs130lp_o41ai_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_o41ai_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.055 3.205 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 2.32 2.725 3.025 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.025 1.875 2.12 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 1.025 1.335 2.12 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.47 0.805 1.435 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3969 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.615 0.935 2.105 ;
        RECT 0.155 1.615 0.935 1.785 ;
        RECT 0.155 0.265 0.445 0.595 ;
        RECT 0.155 0.265 0.325 1.785 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.31 -0.085 2.64 0.485 ;
        RECT 1.335 -0.085 1.665 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.905 1.93 3.075 3.415 ;
        RECT 2.65 1.93 3.075 2.14 ;
        RECT 0.235 1.965 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.985 0.665 3.01 0.835 ;
      RECT 2.82 0.345 3.01 0.835 ;
      RECT 1.92 0.345 2.13 0.835 ;
      RECT 0.985 0.345 1.155 0.835 ;
  END
END scs130lp_o41ai_m

MACRO scs130lp_or2_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2_0 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 0.78 1.365 1.825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.585 2.185 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.955 2.345 2.315 3.025 ;
        RECT 2.055 0.28 2.315 3.025 ;
        RECT 1.62 0.28 2.315 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.195 -0.085 1.45 0.61 ;
        RECT 0.3 -0.085 0.595 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.16 2.345 1.785 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.34 2.41 0.935 2.74 ;
      RECT 0.765 0.28 0.935 2.74 ;
      RECT 0.765 2.005 1.885 2.175 ;
      RECT 1.605 1.505 1.885 2.175 ;
      RECT 0.765 0.28 1.025 0.61 ;
  END
END scs130lp_or2_0

MACRO scs130lp_or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2_1 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.2 1.365 1.515 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.145 0.435 1.515 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 0.255 2.315 3.075 ;
        RECT 1.905 0.255 2.315 1.04 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.405 -0.085 1.735 0.69 ;
        RECT 0.34 -0.085 0.67 0.975 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.16 2.025 1.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.34 1.685 0.67 2.21 ;
      RECT 0.34 1.685 1.875 1.855 ;
      RECT 1.545 1.21 1.875 1.855 ;
      RECT 1.545 0.86 1.715 1.855 ;
      RECT 0.84 0.86 1.715 1.03 ;
      RECT 0.84 0.7 1.1 1.03 ;
  END
END scs130lp_or2_1

MACRO scs130lp_or2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2_2 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 1.15 0.975 1.46 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.79 0.405 1.46 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.645 1.005 1.815 1.925 ;
        RECT 1.545 1.765 1.775 3.075 ;
        RECT 1.585 0.255 1.775 1.14 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.4 0.085 ;
        RECT 1.985 -0.085 2.275 1.095 ;
        RECT 1.945 -0.085 2.275 0.835 ;
        RECT 1.04 -0.085 1.37 0.555 ;
        RECT 0.13 -0.085 0.42 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.4 3.415 ;
        RECT 1.945 2.095 2.275 3.415 ;
        RECT 1.985 1.815 2.275 3.415 ;
        RECT 0.96 1.97 1.375 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.26 1.63 0.47 2.26 ;
      RECT 0.26 1.63 1.375 1.8 ;
      RECT 1.185 0.725 1.375 1.8 ;
      RECT 1.185 1.275 1.475 1.605 ;
      RECT 1.185 0.725 1.415 1.605 ;
      RECT 0.59 0.725 1.415 0.895 ;
      RECT 0.59 0.255 0.87 0.895 ;
  END
END scs130lp_or2_2

MACRO scs130lp_or2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2_4 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.61 1.345 1.02 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.44 1.76 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.54 1.755 3.275 1.945 ;
        RECT 2.855 1.065 3.275 1.945 ;
        RECT 1.53 1.065 3.275 1.245 ;
        RECT 2.39 1.755 2.58 3.075 ;
        RECT 2.39 0.255 2.58 1.245 ;
        RECT 1.54 1.755 1.72 3.075 ;
        RECT 1.53 0.255 1.72 1.245 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.75 -0.085 3.08 0.895 ;
        RECT 1.89 -0.085 2.22 0.895 ;
        RECT 1 -0.085 1.33 0.815 ;
        RECT 0.095 -0.085 0.425 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.75 2.115 3.08 3.415 ;
        RECT 1.89 2.115 2.22 3.415 ;
        RECT 0.96 2.27 1.29 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.095 1.93 0.425 3.075 ;
      RECT 0.095 1.93 1.36 2.1 ;
      RECT 1.19 0.985 1.36 2.1 ;
      RECT 1.19 1.415 2.685 1.585 ;
      RECT 0.61 0.985 1.36 1.175 ;
      RECT 0.61 0.255 0.83 1.175 ;
  END
END scs130lp_or2_4

MACRO scs130lp_or2_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.835 2.15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.455 0.44 1.795 1.78 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2394 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.51 2.43 3.235 2.89 ;
        RECT 2.525 1.18 3.235 2.89 ;
        RECT 2.785 0.55 3.115 1.01 ;
        RECT 2.785 0.55 2.955 2.89 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.965 -0.085 2.295 1.01 ;
        RECT 0.135 -0.085 0.465 1.01 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.72 2.43 2.05 3.415 ;
        RECT 0.315 2.32 0.645 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.115 2.09 1.465 2.78 ;
      RECT 1.115 2.09 2.355 2.26 ;
      RECT 2.025 1.59 2.355 2.26 ;
      RECT 1.115 0.55 1.285 2.78 ;
      RECT 0.955 0.55 1.285 1.01 ;
  END
END scs130lp_or2_lp

MACRO scs130lp_or2_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2_lp2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.905 2.14 1.575 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.18 0.93 2.89 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 0.265 3.235 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.115 -0.085 2.445 0.725 ;
        RECT 0.505 -0.085 0.835 0.725 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.13 2.105 2.46 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.11 1.755 1.44 3.065 ;
      RECT 1.11 1.755 2.725 1.925 ;
      RECT 2.395 1.215 2.725 1.925 ;
      RECT 1.11 0.265 1.28 3.065 ;
      RECT 1.11 0.265 1.655 0.725 ;
  END
END scs130lp_or2_lp2

MACRO scs130lp_or2_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2_m 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.21 1.025 1.405 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.765 0.355 1.435 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.555 0.345 1.765 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 1.92 0.085 ;
        RECT 1.125 -0.085 1.335 0.545 ;
        RECT 0.265 -0.085 0.475 0.545 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 1.92 3.415 ;
        RECT 1.125 2.095 1.335 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.615 1.745 0.945 3.025 ;
      RECT 0.335 1.745 0.945 2.295 ;
      RECT 0.335 1.745 1.375 1.915 ;
      RECT 1.205 0.725 1.375 1.915 ;
      RECT 0.695 0.725 1.375 0.895 ;
      RECT 0.695 0.345 0.905 0.895 ;
  END
END scs130lp_or2_m

MACRO scs130lp_or2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2b_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 2.32 1.785 2.955 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.45 0.775 0.93 1.715 ;
        RECT 0.45 0.775 0.91 1.86 ;
    END
  END BN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.465 1.815 2.795 3.075 ;
        RECT 2.525 0.255 2.795 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.975 -0.085 2.355 1.025 ;
        RECT 1.14 -0.085 1.37 0.62 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.955 1.815 2.295 3.415 ;
        RECT 0.56 2.72 0.805 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.08 1.88 1.38 2.21 ;
      RECT 1.08 1.88 1.73 2.12 ;
      RECT 1.54 0.29 1.73 2.12 ;
      RECT 1.54 1.195 2.355 1.525 ;
      RECT 1.54 0.29 1.77 1.525 ;
      RECT 0.085 2.38 0.39 3.05 ;
      RECT 0.975 2.38 1.305 2.955 ;
      RECT 0.085 2.38 1.305 2.55 ;
      RECT 0.085 0.29 0.28 3.05 ;
      RECT 0.085 0.29 0.97 0.605 ;
  END
END scs130lp_or2b_1

MACRO scs130lp_or2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2b_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 1.415 2.775 1.76 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.875 0.47 1.545 ;
    END
  END BN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.08 0.865 1.445 1.045 ;
        RECT 1.08 0.865 1.41 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.03 -0.085 3.36 0.905 ;
        RECT 1.625 -0.085 1.955 0.355 ;
        RECT 0.59 -0.085 0.935 0.355 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.58 2.27 1.84 3.415 ;
        RECT 0.685 2.055 0.91 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.16 1.715 0.49 2.21 ;
      RECT 0.16 1.715 0.82 1.885 ;
      RECT 0.65 0.525 0.82 1.885 ;
      RECT 2.945 1.075 3.635 1.525 ;
      RECT 2.69 1.075 3.635 1.245 ;
      RECT 2.69 0.525 2.86 1.245 ;
      RECT 0.095 0.525 2.86 0.695 ;
      RECT 0.095 0.29 0.42 0.695 ;
      RECT 2.73 1.93 3.06 2.26 ;
      RECT 1.58 1.93 3.06 2.1 ;
      RECT 1.58 1.155 1.83 2.1 ;
      RECT 1.615 0.865 1.83 2.1 ;
      RECT 1.615 0.865 2.52 1.125 ;
  END
END scs130lp_or2b_2

MACRO scs130lp_or2b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2b_4 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.585 1.425 2.275 1.76 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.295 0.545 2.13 ;
    END
  END BN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.58 1.755 4.235 1.945 ;
        RECT 3.965 1.065 4.235 1.945 ;
        RECT 2.96 1.065 4.235 1.245 ;
        RECT 3.5 1.755 3.69 3.075 ;
        RECT 2.96 0.735 3.69 1.245 ;
        RECT 3.5 0.255 3.69 1.245 ;
        RECT 2.57 0.735 3.69 0.905 ;
        RECT 2.58 1.755 2.83 3.075 ;
        RECT 2.57 0.255 2.83 0.905 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.86 -0.085 4.19 0.895 ;
        RECT 3 -0.085 3.33 0.565 ;
        RECT 2.135 -0.085 2.4 0.905 ;
        RECT 1.24 -0.085 1.57 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.86 2.115 4.19 3.415 ;
        RECT 3 2.115 3.33 3.415 ;
        RECT 2.08 1.93 2.41 3.415 ;
        RECT 0.525 2.64 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.24 1.93 1.57 3.075 ;
      RECT 1.24 1.075 1.415 3.075 ;
      RECT 2.445 1.415 3.795 1.585 ;
      RECT 2.445 1.075 2.79 1.585 ;
      RECT 1.24 1.075 2.79 1.255 ;
      RECT 1.74 0.255 1.965 1.255 ;
      RECT 0.095 2.3 0.355 2.915 ;
      RECT 0.095 2.3 1.045 2.47 ;
      RECT 0.715 0.255 1.045 2.47 ;
  END
END scs130lp_or2b_4

MACRO scs130lp_or2b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2b_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.215 2.555 2.89 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.56 1.175 0.89 1.845 ;
    END
  END BN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.265 2.025 3.715 3.065 ;
        RECT 3.35 0.265 3.715 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.53 -0.085 2.86 0.685 ;
        RECT 0.92 -0.085 1.25 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.735 2.025 3.065 3.415 ;
        RECT 0.66 2.025 0.99 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.43 2.025 1.865 3.065 ;
      RECT 1.695 0.265 1.865 3.065 ;
      RECT 2.835 0.865 3.165 1.535 ;
      RECT 1.695 0.865 3.165 1.035 ;
      RECT 1.695 0.265 2.07 1.035 ;
      RECT 0.13 0.265 0.38 3.065 ;
      RECT 1.185 0.825 1.515 1.495 ;
      RECT 0.13 0.825 1.515 0.995 ;
      RECT 0.13 0.265 0.46 0.995 ;
  END
END scs130lp_or2b_lp

MACRO scs130lp_or2b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or2b_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 2.32 1.765 2.93 ;
    END
  END A
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.21 0.47 2.12 ;
    END
  END BN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.231 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.455 2 2.725 2.86 ;
        RECT 2.535 0.44 2.725 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.945 -0.085 2.275 0.58 ;
        RECT 1.01 -0.085 1.22 0.64 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.945 1.93 2.275 3.415 ;
        RECT 0.525 2.65 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.08 1.93 1.765 2.14 ;
      RECT 1.595 0.47 1.765 2.14 ;
      RECT 2.185 0.86 2.355 1.53 ;
      RECT 1.595 0.86 2.355 1.03 ;
      RECT 1.4 0.47 1.765 0.68 ;
      RECT 0.155 2.3 0.345 2.79 ;
      RECT 0.155 2.3 0.83 2.47 ;
      RECT 0.66 0.5 0.83 2.47 ;
      RECT 1.245 0.86 1.415 1.53 ;
      RECT 0.66 0.86 1.415 1.03 ;
      RECT 0.5 0.5 0.83 0.71 ;
  END
END scs130lp_or2b_m

MACRO scs130lp_or3_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3_0 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.195 1.835 1.865 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 1.135 1.355 1.865 ;
        RECT 1.035 0.805 1.3 1.865 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 0.805 0.865 1.86 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2977 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.42 2.385 2.795 3.065 ;
        RECT 2.545 0.32 2.795 3.065 ;
        RECT 2.33 0.32 2.795 0.65 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.9 -0.085 2.16 0.65 ;
        RECT 0.555 -0.085 1.3 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.665 2.385 2.25 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.5 2.035 0.83 2.78 ;
      RECT 0.105 2.035 0.83 2.34 ;
      RECT 0.105 2.035 2.375 2.215 ;
      RECT 2.015 1.545 2.375 2.215 ;
      RECT 0.105 0.32 0.385 2.34 ;
      RECT 2.015 0.82 2.185 2.215 ;
      RECT 1.47 0.82 2.185 1.005 ;
      RECT 1.47 0.32 1.73 1.005 ;
  END
END scs130lp_or3_0

MACRO scs130lp_or3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3_1 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 1.425 1.895 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.02 1.425 1.33 1.75 ;
        RECT 1.02 0.765 1.295 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.495 0.78 0.845 1.75 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 0.255 2.785 3.075 ;
        RECT 2.38 0.255 2.785 0.905 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.885 -0.085 2.21 0.915 ;
        RECT 0.655 -0.085 1.295 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.66 2.31 2.355 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.92 0.66 2.77 ;
      RECT 0.085 1.92 2.355 2.14 ;
      RECT 2.115 1.085 2.355 2.14 ;
      RECT 0.085 0.28 0.325 2.77 ;
      RECT 1.465 1.085 2.355 1.255 ;
      RECT 1.465 0.28 1.715 1.255 ;
      RECT 0.085 0.28 0.485 0.61 ;
  END
END scs130lp_or3_1

MACRO scs130lp_or3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.515 1.13 1.965 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.045 1.04 1.345 2.12 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.13 0.875 2.12 ;
        RECT 0.425 1.13 0.875 1.775 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.385 1.87 2.725 3.075 ;
        RECT 2.355 0.91 2.685 1.16 ;
        RECT 2.385 0.91 2.64 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.9 -0.085 3.23 0.4 ;
        RECT 1.845 -0.085 2.175 0.4 ;
        RECT 0.565 -0.085 1.235 0.53 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.895 1.815 3.145 3.415 ;
        RECT 1.515 1.92 2.215 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.085 1.945 0.455 2.275 ;
      RECT 0.085 0.345 0.255 2.275 ;
      RECT 2.81 1.33 3.255 1.58 ;
      RECT 2.855 0.57 3.255 1.58 ;
      RECT 0.085 0.7 2.08 0.87 ;
      RECT 1.405 0.57 3.255 0.74 ;
      RECT 0.085 0.345 0.395 0.87 ;
      RECT 1.405 0.28 1.665 0.87 ;
  END
END scs130lp_or3_2

MACRO scs130lp_or3_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3_4 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.345 1.81 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.345 1.355 1.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.375 0.855 1.75 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.32 1.775 4.165 1.945 ;
        RECT 3.985 0.355 4.165 1.945 ;
        RECT 2.32 1.075 4.165 1.245 ;
        RECT 3.98 0.355 4.165 1.245 ;
        RECT 3.18 0.255 3.405 1.245 ;
        RECT 3.18 1.775 3.37 3.075 ;
        RECT 2.32 1.775 2.51 3.075 ;
        RECT 2.32 0.255 2.51 1.245 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.575 -0.085 3.81 0.905 ;
        RECT 2.68 -0.085 3.01 0.905 ;
        RECT 1.765 -0.085 2.13 0.825 ;
        RECT 0.81 -0.085 1.14 0.825 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.54 2.115 3.87 3.415 ;
        RECT 2.68 2.115 3.01 3.415 ;
        RECT 1.745 2.27 2.1 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.345 1.92 0.675 3.075 ;
      RECT 0.345 1.92 2.15 2.1 ;
      RECT 1.98 0.995 2.15 2.1 ;
      RECT 1.98 1.425 3.815 1.595 ;
      RECT 0.345 0.995 2.15 1.165 ;
      RECT 1.31 0.255 1.595 1.165 ;
      RECT 0.345 0.255 0.64 1.165 ;
  END
END scs130lp_or3_4

MACRO scs130lp_or3_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.215 2.275 2.89 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.455 1.215 2.785 2.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.215 3.355 1.885 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.44 0.845 3.065 ;
        RECT 0.125 0.265 0.565 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.605 -0.085 2.935 0.685 ;
        RECT 1.025 -0.085 1.355 0.685 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.045 2.025 1.375 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3.25 2.065 3.725 3.065 ;
      RECT 3.555 0.265 3.725 3.065 ;
      RECT 1.025 0.865 1.355 1.84 ;
      RECT 1.025 0.865 3.725 1.035 ;
      RECT 3.395 0.265 3.725 1.035 ;
      RECT 1.815 0.265 2.145 1.035 ;
  END
END scs130lp_or3_lp

MACRO scs130lp_or3_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3_m 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.075 1.98 1.585 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.765 1.315 1.435 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 0.47 0.805 1.435 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.315 2.155 2.725 2.86 ;
        RECT 2.555 0.275 2.725 2.86 ;
        RECT 2.315 0.275 2.725 0.485 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
      LAYER li ;
        RECT 0 -0.085 2.88 0.085 ;
        RECT 1.905 -0.085 2.115 0.545 ;
        RECT 0.985 -0.085 1.315 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
      LAYER li ;
        RECT 0 3.245 2.88 3.415 ;
        RECT 1.805 2.155 2.135 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.295 1.795 1.625 3.025 ;
      RECT 0.685 1.795 0.895 2.295 ;
      RECT 0.235 1.795 2.33 1.965 ;
      RECT 2.16 0.725 2.33 1.965 ;
      RECT 0.235 0.345 0.425 1.965 ;
      RECT 1.495 0.725 2.33 0.895 ;
      RECT 1.495 0.345 1.685 0.895 ;
  END
END scs130lp_or3_m

MACRO scs130lp_or3b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3b_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.43 2.64 2.325 3.02 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 0.84 1.975 2.13 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.405 2.49 ;
    END
  END CN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.975 1.815 3.255 3.075 ;
        RECT 3.085 0.35 3.255 3.075 ;
        RECT 2.975 0.35 3.255 1.16 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.495 -0.085 2.755 1.15 ;
        RECT 1.56 -0.085 1.79 0.67 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.495 1.82 2.755 3.415 ;
        RECT 0.095 2.66 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.06 2.3 2.325 2.47 ;
      RECT 2.155 0.39 2.325 2.47 ;
      RECT 1.06 1.88 1.39 2.47 ;
      RECT 1.22 0.42 1.39 2.47 ;
      RECT 2.155 1.32 2.905 1.65 ;
      RECT 1.06 0.42 1.39 0.75 ;
      RECT 1.96 0.39 2.325 0.67 ;
      RECT 0.595 0.395 0.855 2.935 ;
      RECT 0.595 1 1.05 1.67 ;
  END
END scs130lp_or3b_1

MACRO scs130lp_or3b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3b_2 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.91 1.425 2.305 2.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 1.125 2.815 2.12 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.405 0.58 1.75 ;
    END
  END CN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.1 1.815 1.575 2.12 ;
        RECT 1.1 0.255 1.36 1.01 ;
        RECT 1.1 0.255 1.27 2.12 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.485 -0.085 2.815 0.615 ;
        RECT 1.53 -0.085 1.93 0.895 ;
        RECT 0.555 -0.085 0.93 0.895 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.675 2.64 2.005 3.415 ;
        RECT 0.815 2.64 1.145 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.985 0.28 3.265 2.3 ;
      RECT 1.44 1.19 1.72 1.52 ;
      RECT 2.1 0.28 2.305 1.235 ;
      RECT 1.55 1.065 2.305 1.235 ;
      RECT 2.1 0.785 3.265 0.955 ;
      RECT 2.1 0.28 2.315 0.955 ;
      RECT 2.485 2.29 2.815 2.965 ;
      RECT 0.29 2.29 2.815 2.46 ;
      RECT 0.29 1.92 0.93 2.46 ;
      RECT 0.75 1.065 0.93 2.46 ;
      RECT 0.125 1.065 0.93 1.235 ;
      RECT 0.125 0.7 0.385 1.235 ;
  END
END scs130lp_or3b_2

MACRO scs130lp_or3b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3b_4 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.02 1.345 3.275 2.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.445 1.345 3.74 2.145 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 0.47 0.835 2.12 ;
    END
  END CN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.005 1.815 2.725 2.145 ;
        RECT 1.005 1.075 2.51 1.245 ;
        RECT 2.32 0.255 2.51 1.245 ;
        RECT 1.43 0.255 1.65 1.245 ;
        RECT 1.005 1.075 1.185 2.145 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.675 -0.085 4.005 0.835 ;
        RECT 2.72 -0.085 3.05 0.835 ;
        RECT 1.82 -0.085 2.15 0.905 ;
        RECT 1.005 -0.085 1.26 0.905 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 2.77 2.655 3.1 3.415 ;
        RECT 1.855 2.655 2.185 3.415 ;
        RECT 0.995 2.655 1.325 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.155 2.76 4.71 3.075 ;
      RECT 4.53 0.255 4.71 3.075 ;
      RECT 4.26 1.815 4.71 3.075 ;
      RECT 1.355 1.415 2.85 1.645 ;
      RECT 2.68 1.005 2.85 1.645 ;
      RECT 2.68 1.005 4.71 1.175 ;
      RECT 4.175 0.255 4.71 1.175 ;
      RECT 3.22 0.255 3.505 1.175 ;
      RECT 0.205 2.315 4.09 2.485 ;
      RECT 3.92 1.345 4.09 2.485 ;
      RECT 0.205 0.71 0.455 2.485 ;
      RECT 3.92 1.345 4.36 1.645 ;
  END
END scs130lp_or3b_4

MACRO scs130lp_or3b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3b_lp 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.035 3.715 1.41 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.81 1.675 3.715 2.15 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.445 1.175 0.835 1.845 ;
    END
  END CN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.445 0.44 4.685 2.89 ;
        RECT 4.245 2.075 4.575 3.065 ;
        RECT 4.355 0.44 4.685 0.945 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.565 -0.085 3.895 0.855 ;
        RECT 1.875 0.895 2.405 1.145 ;
        RECT 2.235 -0.085 2.405 1.145 ;
        RECT 0.905 -0.085 1.235 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.605 2.68 3.935 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.825 1.325 2.155 2.715 ;
      RECT 2.46 2.33 4.065 2.5 ;
      RECT 3.895 1.225 4.065 2.5 ;
      RECT 2.46 1.325 2.63 2.5 ;
      RECT 3.895 1.225 4.225 1.895 ;
      RECT 1.525 1.325 2.825 1.495 ;
      RECT 2.655 0.485 2.825 1.495 ;
      RECT 1.525 0.265 1.695 1.495 ;
      RECT 2.655 0.485 3.075 0.855 ;
      RECT 1.525 0.265 2.055 0.675 ;
      RECT 1.295 2.895 2.915 3.065 ;
      RECT 2.585 2.68 2.915 3.065 ;
      RECT 1.295 1.845 1.625 3.065 ;
      RECT 0.095 2.025 0.445 3.065 ;
      RECT 0.095 0.265 0.265 3.065 ;
      RECT 1.015 0.825 1.345 1.45 ;
      RECT 0.095 0.825 1.345 0.995 ;
      RECT 0.095 0.265 0.445 0.995 ;
  END
END scs130lp_or3b_lp

MACRO scs130lp_or3b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or3b_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 2.67 2.345 3 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.21 2.035 1.75 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.49 ;
    END
  END CN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.231 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.925 2.2 3.205 2.86 ;
        RECT 3.035 0.265 3.205 2.86 ;
        RECT 2.86 0.265 3.205 0.595 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.43 -0.085 2.64 0.55 ;
        RECT 1.57 -0.085 1.78 0.55 ;
        RECT 0.165 -0.085 0.375 0.585 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.53 2.28 2.7 3.415 ;
        RECT 2.37 2.28 2.7 2.49 ;
        RECT 0.165 2.785 0.355 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.02 2.13 1.7 2.34 ;
      RECT 1.53 1.93 1.7 2.34 ;
      RECT 1.18 0.35 1.35 2.34 ;
      RECT 1.53 1.93 2.745 2.1 ;
      RECT 2.575 0.775 2.745 2.1 ;
      RECT 2.575 0.775 2.855 1.445 ;
      RECT 2 0.775 2.855 0.945 ;
      RECT 2 0.37 2.21 0.945 ;
      RECT 1.14 0.35 1.35 0.68 ;
      RECT 0.595 0.385 0.805 2.985 ;
      RECT 0.595 1.23 0.925 1.9 ;
  END
END scs130lp_or3b_m

MACRO scs130lp_or4_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 1.2 2.285 1.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.12 1.83 1.485 ;
        RECT 1.465 0.805 1.805 1.485 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 1.57 1.295 2.22 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.805 0.365 2.13 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2998 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.775 2.39 3.275 3.075 ;
        RECT 3.025 0.305 3.275 3.075 ;
        RECT 2.76 0.305 3.275 0.635 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.315 -0.085 2.59 0.635 ;
        RECT 1.08 -0.085 1.665 0.635 ;
        RECT 0.17 -0.085 0.47 0.635 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.92 2.39 2.605 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.2 2.455 1.635 2.785 ;
      RECT 1.465 2.05 1.635 2.785 ;
      RECT 0.535 2.43 1.635 2.785 ;
      RECT 0.535 1.23 0.705 2.785 ;
      RECT 1.465 2.05 2.76 2.22 ;
      RECT 2.465 0.86 2.76 2.22 ;
      RECT 2.465 0.86 2.855 1.53 ;
      RECT 0.64 0.305 0.9 1.4 ;
      RECT 1.975 0.86 2.855 1.03 ;
      RECT 1.975 0.305 2.145 1.03 ;
      RECT 1.835 0.305 2.145 0.635 ;
  END
END scs130lp_or4_0

MACRO scs130lp_or4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.995 1.425 2.325 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.395 1.005 1.775 1.83 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.585 0.985 1.155 1.83 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.78 0.41 1.83 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 0.255 3.275 3.075 ;
        RECT 2.7 0.255 3.275 0.905 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.285 -0.085 2.53 0.905 ;
        RECT 0.99 -0.085 1.66 0.475 ;
        RECT 0.13 -0.085 0.43 0.61 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.67 2.445 2.835 3.415 ;
        RECT 2.505 2.32 2.835 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.16 2 0.49 2.775 ;
      RECT 0.16 2 2.335 2.26 ;
      RECT 2.565 1.075 2.815 2.15 ;
      RECT 2.165 1.93 2.815 2.15 ;
      RECT 1.945 1.075 2.815 1.245 ;
      RECT 1.945 0.28 2.115 1.245 ;
      RECT 0.6 0.645 2.115 0.815 ;
      RECT 1.83 0.28 2.115 0.815 ;
      RECT 0.6 0.28 0.82 0.815 ;
  END
END scs130lp_or4_1

MACRO scs130lp_or4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.005 1.355 2.395 1.675 ;
        RECT 2.005 2.345 2.355 2.96 ;
        RECT 2.005 1.355 2.245 2.96 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.52 1.005 1.835 2.96 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 1.075 1.35 2.96 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.76 0.365 1.75 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5943 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 1.105 3.26 3.075 ;
        RECT 3.03 0.255 3.26 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.43 -0.085 3.72 1.105 ;
        RECT 2.455 -0.085 2.86 0.845 ;
        RECT 2.19 -0.085 2.86 0.485 ;
        RECT 1.26 -0.085 1.59 0.485 ;
        RECT 0.3 -0.085 0.63 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.43 1.815 3.72 3.415 ;
        RECT 2.525 1.845 2.855 3.415 ;
        RECT 2.415 1.845 2.855 2.175 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.32 1.92 0.705 2.21 ;
      RECT 0.535 0.735 0.705 2.21 ;
      RECT 2.575 1.285 2.855 1.615 ;
      RECT 2.575 1.015 2.745 1.615 ;
      RECT 2.005 1.015 2.745 1.185 ;
      RECT 2.005 0.655 2.285 1.185 ;
      RECT 0.535 0.735 0.98 0.905 ;
      RECT 1.76 0.255 2.02 0.825 ;
      RECT 0.8 0.655 2.285 0.825 ;
      RECT 0.8 0.255 1.09 0.825 ;
  END
END scs130lp_or4_2

MACRO scs130lp_or4_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4_4 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2 1.345 2.255 1.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 1.345 1.83 1.76 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.425 1.325 1.76 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.455 1.76 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.765 1.765 4.715 1.935 ;
        RECT 4.455 0.47 4.715 1.935 ;
        RECT 4.43 1.085 4.715 1.935 ;
        RECT 2.765 1.085 4.715 1.255 ;
        RECT 3.625 0.255 3.85 1.255 ;
        RECT 3.625 1.765 3.815 3.075 ;
        RECT 2.765 1.765 2.955 3.075 ;
        RECT 2.765 0.255 2.955 1.255 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 4.02 -0.085 4.285 0.915 ;
        RECT 3.125 -0.085 3.455 0.915 ;
        RECT 2.19 -0.085 2.52 0.825 ;
        RECT 1.19 -0.085 1.52 0.825 ;
        RECT 0.25 -0.085 0.58 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.985 2.105 4.315 3.415 ;
        RECT 3.125 2.105 3.455 3.415 ;
        RECT 2.185 2.27 2.515 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.25 1.93 0.58 3.075 ;
      RECT 0.25 1.93 2.595 2.1 ;
      RECT 2.425 0.995 2.595 2.1 ;
      RECT 2.425 1.425 4.26 1.595 ;
      RECT 0.75 0.995 2.595 1.165 ;
      RECT 1.69 0.255 2.02 1.165 ;
      RECT 0.75 0.255 1.01 1.165 ;
  END
END scs130lp_or4_4

MACRO scs130lp_or4_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4_lp 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.675 3.37 2.89 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.675 2.275 2.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.01 1.265 1.34 2.89 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.44 1.205 0.83 1.875 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.355 0.44 4.685 2.89 ;
        RECT 4.08 2.075 4.41 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.565 -0.085 3.895 1.145 ;
        RECT 1.87 0.895 2.455 1.145 ;
        RECT 2.285 -0.085 2.455 1.145 ;
        RECT 0.905 -0.085 1.235 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.55 2.075 3.88 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.09 2.075 0.545 3.065 ;
      RECT 0.09 0.265 0.26 3.065 ;
      RECT 3.845 1.325 4.175 1.695 ;
      RECT 1.52 1.325 4.175 1.495 ;
      RECT 2.775 0.815 3.105 1.495 ;
      RECT 1.52 0.265 1.69 1.495 ;
      RECT 0.09 0.855 1.69 1.025 ;
      RECT 1.52 0.265 2.105 0.675 ;
      RECT 0.09 0.265 0.445 0.675 ;
  END
END scs130lp_or4_lp

MACRO scs130lp_or4_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1 2.46 1.51 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 0.84 1.895 1.38 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 0.47 1.285 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 0.84 0.355 2.49 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.795 2.155 3.265 2.86 ;
        RECT 3.035 0.28 3.265 2.86 ;
        RECT 2.935 0.28 3.265 0.47 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.425 -0.085 2.755 0.465 ;
        RECT 1.465 -0.085 1.795 0.485 ;
        RECT 0.225 -0.085 0.555 0.485 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.285 2.155 2.615 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.775 1.795 2.105 3.025 ;
      RECT 0.6 1.965 0.905 2.295 ;
      RECT 2.64 0.65 2.81 1.965 ;
      RECT 0.735 1.795 2.81 1.965 ;
      RECT 0.735 0.345 0.925 1.965 ;
      RECT 2.075 0.65 2.81 0.82 ;
      RECT 1.975 0.33 2.245 0.66 ;
  END
END scs130lp_or4_m

MACRO scs130lp_or4b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4b_1 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 1.85 2.735 2.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.295 2.725 0.655 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.725 1.58 2.305 3.075 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.555 0.48 2.235 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.335 1.815 3.755 3.075 ;
        RECT 3.485 0.255 3.755 3.075 ;
        RECT 3.405 0.255 3.755 1.095 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.895 -0.085 3.235 1.07 ;
        RECT 1.705 -0.085 1.905 1.03 ;
        RECT 0.78 -0.085 1.01 1.03 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.905 1.815 3.165 3.415 ;
        RECT 0.745 2.745 1.04 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.06 1.88 1.545 2.21 ;
      RECT 1.365 1.24 1.545 2.21 ;
      RECT 2.96 1.24 3.315 1.625 ;
      RECT 1.365 1.24 3.315 1.41 ;
      RECT 2.32 0.825 2.65 1.41 ;
      RECT 1.365 0.7 1.535 2.21 ;
      RECT 1.18 0.7 1.535 1.03 ;
      RECT 0.28 2.405 0.575 3.03 ;
      RECT 0.28 2.405 0.89 2.575 ;
      RECT 0.65 1.215 0.89 2.575 ;
      RECT 0.65 1.215 1.195 1.545 ;
      RECT 0.28 1.215 1.195 1.385 ;
      RECT 0.28 0.7 0.61 1.385 ;
  END
END scs130lp_or4b_1

MACRO scs130lp_or4b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4b_2 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.85 1.345 2.275 1.835 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.445 0.84 2.765 1.835 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 1.125 3.245 1.835 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.375 0.48 1.75 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.14 0.255 1.33 1.155 ;
        RECT 1.01 1.845 1.32 2.185 ;
        RECT 1.01 0.985 1.18 2.185 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.485 -0.085 3.745 0.555 ;
        RECT 2.455 -0.085 2.815 0.61 ;
        RECT 1.5 -0.085 1.89 0.835 ;
        RECT 0.64 -0.085 0.97 0.815 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 1.5 2.695 1.83 3.415 ;
        RECT 0.64 2.695 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.5 2.005 3.745 2.185 ;
      RECT 3.415 0.725 3.745 2.185 ;
      RECT 1.5 1.005 1.67 2.185 ;
      RECT 1.35 1.335 1.67 1.665 ;
      RECT 1.5 1.005 2.275 1.175 ;
      RECT 2.06 0.28 2.275 1.175 ;
      RECT 2.985 0.725 3.745 0.895 ;
      RECT 2.985 0.255 3.315 0.895 ;
      RECT 3.1 2.355 3.44 3.045 ;
      RECT 0.66 2.355 3.44 2.525 ;
      RECT 0.66 0.985 0.83 2.525 ;
      RECT 0.115 1.92 0.83 2.26 ;
      RECT 0.65 0.985 0.83 2.26 ;
      RECT 0.115 0.985 0.83 1.155 ;
      RECT 0.115 0.7 0.445 1.155 ;
  END
END scs130lp_or4b_2

MACRO scs130lp_or4b_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4b_4 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.345 2.315 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.385 1.92 2.855 2.94 ;
        RECT 2.485 1.345 2.855 2.94 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 1.345 3.685 2.94 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.73 1.535 5.195 2.205 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.47 1.695 1.715 3.075 ;
        RECT 0.61 0.655 1.68 0.825 ;
        RECT 1.47 0.485 1.68 0.825 ;
        RECT 0.09 1.695 1.715 1.865 ;
        RECT 0.61 1.695 0.8 3.075 ;
        RECT 0.61 0.255 0.8 0.825 ;
        RECT 0.09 1.005 0.79 1.175 ;
        RECT 0.61 0.255 0.79 1.175 ;
        RECT 0.09 1.005 0.335 1.865 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.205 -0.085 4.7 1.015 ;
        RECT 3.93 -0.085 4.7 0.835 ;
        RECT 2.73 -0.085 3.4 0.825 ;
        RECT 1.85 -0.085 2.18 0.825 ;
        RECT 0.97 -0.085 1.3 0.485 ;
        RECT 0.11 -0.085 0.44 0.835 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 4.425 2.715 4.755 3.415 ;
        RECT 1.885 1.92 2.215 3.415 ;
        RECT 0.97 2.035 1.3 3.415 ;
        RECT 0.11 2.035 0.44 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 4.925 2.375 5.185 3.075 ;
      RECT 4.26 2.375 5.185 2.545 ;
      RECT 4.26 1.185 4.56 2.545 ;
      RECT 4.215 1.185 4.56 1.515 ;
      RECT 4.215 1.185 5.13 1.355 ;
      RECT 4.87 0.7 5.13 1.355 ;
      RECT 3.855 1.815 4.09 3.075 ;
      RECT 3.855 1.005 4.035 3.075 ;
      RECT 0.505 1.355 1.905 1.525 ;
      RECT 1.735 0.995 1.905 1.525 ;
      RECT 1.735 1.005 4.035 1.175 ;
      RECT 1.735 0.995 3.76 1.175 ;
      RECT 3.57 0.255 3.76 1.175 ;
      RECT 2.35 0.255 2.56 1.175 ;
  END
END scs130lp_or4b_4

MACRO scs130lp_or4b_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4b_lp 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 1.255 4.195 1.925 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.935 1.255 3.265 2.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.255 2.755 2.89 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.455 1.175 0.835 1.845 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4005 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.375 2.065 5.175 3.065 ;
        RECT 4.925 0.265 5.175 3.065 ;
        RECT 4.845 0.265 5.175 0.725 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
      LAYER li ;
        RECT 0 -0.085 5.28 0.085 ;
        RECT 4.055 -0.085 4.385 0.725 ;
        RECT 2.475 -0.085 2.805 0.725 ;
        RECT 0.895 -0.085 1.225 0.645 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
      LAYER li ;
        RECT 0 3.245 5.28 3.415 ;
        RECT 3.755 2.105 4.085 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.535 2.065 1.865 3.065 ;
      RECT 1.685 0.265 1.865 3.065 ;
      RECT 4.375 0.905 4.705 1.84 ;
      RECT 1.685 0.905 4.705 1.075 ;
      RECT 3.265 0.265 3.595 1.075 ;
      RECT 1.685 0.265 2.015 1.075 ;
      RECT 0.105 2.025 0.445 3.065 ;
      RECT 0.105 0.265 0.275 3.065 ;
      RECT 1.175 0.825 1.505 1.495 ;
      RECT 0.105 0.825 1.505 0.995 ;
      RECT 0.105 0.265 0.435 0.995 ;
  END
END scs130lp_or4b_lp

MACRO scs130lp_or4b_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4b_m 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 1.575 3.205 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 0.265 2.725 0.64 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 2.69 2.245 3.025 ;
    END
  END C
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.49 0.47 2.16 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.345 1.93 3.685 2.86 ;
        RECT 3.385 0.47 3.685 2.86 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 2.905 -0.085 3.115 0.935 ;
        RECT 1.595 -0.085 1.805 0.935 ;
        RECT 0.66 -0.085 0.87 0.935 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 2.995 2.155 3.165 3.415 ;
        RECT 2.835 2.155 3.165 2.365 ;
        RECT 0.58 2.69 0.91 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.485 2.855 2.815 3.025 ;
      RECT 2.485 2.005 2.655 3.025 ;
      RECT 1.245 2.005 2.655 2.335 ;
      RECT 1.245 0.75 1.415 2.335 ;
      RECT 1.245 1.225 2.715 1.395 ;
      RECT 2.385 0.835 2.715 1.395 ;
      RECT 1.05 0.75 1.415 0.96 ;
      RECT 0.21 2.34 0.4 2.83 ;
      RECT 0.21 2.34 0.82 2.51 ;
      RECT 0.65 1.14 0.82 2.51 ;
      RECT 0.65 1.14 1.065 1.825 ;
      RECT 0.15 1.14 1.065 1.31 ;
      RECT 0.15 0.795 0.48 1.31 ;
  END
END scs130lp_or4b_m

MACRO scs130lp_or4bb_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4bb_1 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.06 2.305 3.205 2.995 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.475 0.78 2.975 1.025 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.435 0.765 0.92 1.435 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.56 2.045 1.335 2.55 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.895 1.815 4.235 3.075 ;
        RECT 3.965 0.255 4.235 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.495 -0.085 3.795 1.025 ;
        RECT 2.43 -0.085 2.76 0.61 ;
        RECT 1.55 -0.085 1.86 0.605 ;
        RECT 0.67 -0.085 0.92 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.375 1.815 3.675 3.415 ;
        RECT 0.56 2.72 0.82 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.62 1.965 1.89 2.33 ;
      RECT 1.62 1.965 2.965 2.135 ;
      RECT 2.795 1.195 2.965 2.135 ;
      RECT 2.795 1.195 3.795 1.525 ;
      RECT 2.03 1.195 3.795 1.365 ;
      RECT 3.155 0.28 3.325 1.525 ;
      RECT 2.03 0.28 2.26 1.365 ;
      RECT 2.94 0.28 3.325 0.61 ;
      RECT 0.085 1.615 0.39 3.05 ;
      RECT 0.085 1.615 2.615 1.795 ;
      RECT 2.285 1.535 2.615 1.795 ;
      RECT 0.085 0.28 0.265 3.05 ;
      RECT 0.085 0.28 0.5 0.595 ;
      RECT 1.53 0.775 1.86 1.435 ;
      RECT 1.09 0.775 1.86 0.945 ;
      RECT 1.09 0.28 1.36 0.945 ;
      RECT 0.99 2.72 1.785 3.05 ;
  END
END scs130lp_or4bb_1

MACRO scs130lp_or4bb_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4bb_2 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.035 0.775 1.31 1.445 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.5 0.925 1.92 1.455 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.58 0.47 0.815 1.435 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.215 1.405 4.715 1.76 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.45 0.255 3.695 2.275 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.8 0.085 ;
        RECT 3.865 -0.085 4.14 0.895 ;
        RECT 2.98 -0.085 3.28 1.015 ;
        RECT 1.865 -0.085 2.195 0.415 ;
        RECT 0.985 -0.085 1.245 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.8 3.415 ;
        RECT 3.845 2.785 4.175 3.415 ;
        RECT 2.985 2.785 3.315 3.415 ;
        RECT 0.96 2.045 1.255 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.475 2.445 2.805 3.075 ;
      RECT 2.475 2.445 4.205 2.615 ;
      RECT 3.865 1.93 4.205 2.615 ;
      RECT 3.865 1.93 4.7 2.26 ;
      RECT 3.865 1.065 4.035 2.615 ;
      RECT 3.865 1.065 4.665 1.235 ;
      RECT 4.335 0.7 4.665 1.235 ;
      RECT 2.435 1.995 2.81 2.275 ;
      RECT 2.64 0.28 2.81 2.275 ;
      RECT 2.64 1.185 3.28 1.515 ;
      RECT 1.48 0.585 2.81 0.755 ;
      RECT 2.435 0.28 2.81 0.755 ;
      RECT 1.415 0.265 1.65 0.595 ;
      RECT 0.495 1.625 0.79 2.39 ;
      RECT 0.16 1.625 2.46 1.795 ;
      RECT 2.13 0.925 2.46 1.795 ;
      RECT 0.16 0.28 0.41 1.795 ;
  END
END scs130lp_or4bb_2

MACRO scs130lp_or4bb_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4bb_4 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.02 1.21 1.355 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.525 1.345 1.89 1.755 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.21 0.365 1.75 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.875 0.955 6.155 1.75 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.79 1.745 5.225 1.915 ;
        RECT 4.89 0.895 5.225 1.915 ;
        RECT 3.465 0.895 5.225 1.145 ;
        RECT 4.65 1.745 4.84 3.075 ;
        RECT 3.79 1.745 3.98 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 4.99 -0.085 5.32 0.385 ;
        RECT 3.955 -0.085 4.285 0.385 ;
        RECT 2.88 -0.085 3.21 0.385 ;
        RECT 1.865 -0.085 2.195 0.815 ;
        RECT 0.875 -0.085 1.195 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.01 2.085 5.34 3.415 ;
        RECT 4.15 2.085 4.48 3.415 ;
        RECT 3.29 2.095 3.62 3.415 ;
        RECT 0.895 2.265 1.225 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 5.51 1.92 5.865 2.21 ;
      RECT 5.51 0.555 5.705 2.21 ;
      RECT 2.87 0.555 3.13 1.545 ;
      RECT 2.87 0.555 5.705 0.725 ;
      RECT 5.535 0.31 5.865 0.715 ;
      RECT 2.765 1.755 3.095 3.075 ;
      RECT 2.53 1.755 3.54 1.925 ;
      RECT 3.3 1.325 3.54 1.925 ;
      RECT 2.53 0.255 2.7 1.925 ;
      RECT 3.3 1.325 4.72 1.575 ;
      RECT 1.525 0.995 2.7 1.165 ;
      RECT 2.365 0.255 2.7 1.165 ;
      RECT 1.365 0.255 1.695 1.04 ;
      RECT 0.355 1.92 0.685 2.21 ;
      RECT 0.355 1.925 2.35 2.095 ;
      RECT 2.1 1.345 2.35 2.095 ;
      RECT 0.535 0.73 0.705 2.095 ;
      RECT 0.355 0.73 0.705 1.04 ;
  END
END scs130lp_or4bb_4

MACRO scs130lp_or4bb_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4bb_lp 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.405 1.545 5.865 1.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.355 1.815 4.685 2.15 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.4 1.475 1.795 1.805 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.395 1.11 6.725 1.78 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 2.325 0.835 3.065 ;
        RECT 0.125 0.265 0.455 0.595 ;
        RECT 0.125 0.265 0.325 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.2 0.085 ;
        RECT 5.965 -0.085 6.295 0.675 ;
        RECT 5.32 -0.085 5.65 1.365 ;
        RECT 3.66 -0.085 3.99 0.935 ;
        RECT 0.915 -0.085 1.245 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.2 3.415 ;
        RECT 5.845 2.755 6.175 3.415 ;
        RECT 1.035 2.335 1.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.395 2.075 6.725 3.065 ;
      RECT 4.355 2.355 4.685 2.685 ;
      RECT 4.355 2.405 6.725 2.575 ;
      RECT 6.395 2.075 7.085 2.245 ;
      RECT 6.915 0.265 7.085 2.245 ;
      RECT 6.755 0.265 7.085 0.675 ;
      RECT 2.545 2.41 4.175 2.58 ;
      RECT 4.005 1.465 4.175 2.58 ;
      RECT 2.545 1.465 2.715 2.58 ;
      RECT 4.865 2.055 6.215 2.225 ;
      RECT 6.045 0.905 6.215 2.225 ;
      RECT 4.865 1.465 5.035 2.225 ;
      RECT 4.005 1.465 5.035 1.635 ;
      RECT 2.36 1.125 2.69 1.635 ;
      RECT 5.83 0.905 6.215 1.365 ;
      RECT 2.505 2.865 5.155 3.035 ;
      RECT 2.505 2.76 2.835 3.035 ;
      RECT 3.495 1.115 3.825 2.23 ;
      RECT 0.855 1.125 1.13 1.795 ;
      RECT 0.855 1.125 1.945 1.295 ;
      RECT 1.775 0.775 1.945 1.295 ;
      RECT 2.87 1.115 4.34 1.285 ;
      RECT 4.17 0.895 4.34 1.285 ;
      RECT 2.87 0.605 3.2 1.285 ;
      RECT 4.17 0.895 4.78 1.065 ;
      RECT 4.45 0.605 4.78 1.065 ;
      RECT 1.775 0.775 3.2 0.945 ;
      RECT 1.565 1.985 1.895 3.065 ;
      RECT 1.565 1.985 2.365 2.485 ;
      RECT 2.035 1.815 2.365 2.485 ;
      RECT 1.05 1.985 2.365 2.155 ;
      RECT 0.505 1.975 1.22 2.145 ;
      RECT 0.505 0.775 0.675 2.145 ;
      RECT 0.505 0.775 1.595 0.945 ;
      RECT 1.425 0.265 1.595 0.945 ;
      RECT 1.425 0.265 2.035 0.595 ;
  END
END scs130lp_or4bb_lp

MACRO scs130lp_or4bb_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_or4bb_m 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.035 2.015 3.505 2.32 ;
        RECT 3.035 2.015 3.205 2.91 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 0.975 3.015 1.485 ;
    END
  END B
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.455 0.775 0.805 1.445 ;
    END
  END CN
  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.585 2.005 1.16 2.525 ;
    END
  END DN
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2226 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.935 2.32 4.225 2.91 ;
        RECT 4.055 0.345 4.225 2.91 ;
        RECT 3.955 0.345 4.225 0.675 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 4.32 0.085 ;
        RECT 3.545 -0.085 3.735 0.545 ;
        RECT 2.47 -0.085 2.8 0.445 ;
        RECT 1.65 -0.085 1.86 0.545 ;
        RECT 0.7 -0.085 0.91 0.555 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 4.32 3.415 ;
        RECT 3.385 2.595 3.715 3.415 ;
        RECT 0.585 2.76 0.775 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.7 2.175 2.855 2.505 ;
      RECT 2.685 1.665 2.855 2.505 ;
      RECT 2.685 1.665 3.875 1.835 ;
      RECT 3.705 1.025 3.875 1.835 ;
      RECT 3.195 0.345 3.365 1.835 ;
      RECT 2.08 0.625 3.365 0.795 ;
      RECT 3.02 0.345 3.365 0.795 ;
      RECT 2.08 0.365 2.29 0.795 ;
      RECT 0.105 1.625 0.365 2.96 ;
      RECT 0.105 1.625 2.375 1.795 ;
      RECT 2.205 1.365 2.375 1.795 ;
      RECT 0.105 0.265 0.275 2.96 ;
      RECT 0.105 0.265 0.48 0.595 ;
      RECT 1.535 0.735 1.705 1.445 ;
      RECT 1.13 0.735 1.705 0.905 ;
      RECT 1.13 0.355 1.34 0.905 ;
      RECT 1.015 2.695 1.735 3.025 ;
  END
END scs130lp_or4bb_m

MACRO scs130lp_sdfbbn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfbbn_1 0 0 ;
  SIZE 17.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.86 0.87 4.195 1.54 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.49 0.81 1.82 1.82 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 17.315 1.815 17.67 3.065 ;
        RECT 17.5 0.265 17.67 3.065 ;
        RECT 17.315 0.265 17.67 1.125 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5922 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.9 1.835 16.255 3.065 ;
        RECT 16.085 0.265 16.255 3.065 ;
        RECT 15.85 0.265 16.255 1.145 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.005 1.345 15.365 1.78 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.215 0.55 1.885 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.85 1.215 1.31 1.78 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 0.891892 LAYER li ;
      ANTENNAMAXAREACAR 0.891892 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.837838 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.837838 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 13.055 1.18 13.345 1.41 ;
        RECT 8.735 1.225 13.345 1.365 ;
        RECT 8.735 1.18 9.025 1.41 ;
      LAYER li ;
        RECT 13 1.18 13.33 1.78 ;
        RECT 8.57 1.08 8.995 1.41 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.76 0.245 ;
      LAYER li ;
        RECT 0 -0.085 17.76 0.085 ;
        RECT 16.84 -0.085 17.09 0.725 ;
        RECT 15.42 -0.085 15.67 1.145 ;
        RECT 12.645 -0.085 12.975 0.65 ;
        RECT 10.615 -0.085 10.865 0.905 ;
        RECT 7.875 -0.085 8.205 0.525 ;
        RECT 5.465 -0.085 5.795 0.77 ;
        RECT 3.655 -0.085 3.985 0.69 ;
        RECT 2.35 -0.085 2.68 0.995 ;
        RECT 0.155 -0.085 0.485 1.035 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.76 3.575 ;
      LAYER li ;
        RECT 0 3.245 17.76 3.415 ;
        RECT 16.885 1.815 17.135 3.415 ;
        RECT 15.39 2.82 15.72 3.415 ;
        RECT 14.325 2.82 14.655 3.415 ;
        RECT 13.105 2.47 13.355 3.415 ;
        RECT 10.345 1.905 10.675 3.415 ;
        RECT 8.3 2.29 8.63 3.415 ;
        RECT 5.47 2.675 5.8 3.415 ;
        RECT 3.795 2.07 3.965 3.415 ;
        RECT 2.395 2.035 2.565 3.415 ;
        RECT 0.545 2.415 0.795 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 16.455 1.305 16.705 2.495 ;
      RECT 16.455 1.305 17.32 1.635 ;
      RECT 16.455 0.265 16.66 2.495 ;
      RECT 13.535 1.96 13.865 3.065 ;
      RECT 13.535 2.47 15.72 2.64 ;
      RECT 15.55 1.325 15.72 2.64 ;
      RECT 14.05 1.085 14.22 2.64 ;
      RECT 12.64 1.96 13.865 2.29 ;
      RECT 15.55 1.325 15.905 1.655 ;
      RECT 13.905 0.615 14.155 1.255 ;
      RECT 14.4 1.96 15.21 2.29 ;
      RECT 14.4 0.995 14.73 2.29 ;
      RECT 14.4 0.995 15.24 1.165 ;
      RECT 14.91 0.265 15.24 1.165 ;
      RECT 14.335 0.265 14.665 0.815 ;
      RECT 13.235 0.265 13.565 0.65 ;
      RECT 13.235 0.265 14.665 0.435 ;
      RECT 11.47 2.12 11.88 2.715 ;
      RECT 11.71 0.575 11.88 2.715 ;
      RECT 13.54 1.435 13.87 1.765 ;
      RECT 13.54 0.83 13.71 1.765 ;
      RECT 11.47 0.575 11.88 1.165 ;
      RECT 11.47 0.83 13.71 1 ;
      RECT 11.12 2.895 12.43 3.065 ;
      RECT 12.1 1.7 12.43 3.065 ;
      RECT 11.12 1.085 11.29 3.065 ;
      RECT 11.12 1.345 11.53 1.675 ;
      RECT 7.045 0.705 7.31 1.38 ;
      RECT 10.265 1.085 11.29 1.255 ;
      RECT 10.265 0.265 10.435 1.255 ;
      RECT 7.045 0.705 8.555 0.875 ;
      RECT 8.385 0.265 8.555 0.875 ;
      RECT 8.385 0.265 10.435 0.435 ;
      RECT 9.525 1.915 9.855 2.755 ;
      RECT 9.685 1.055 9.855 2.755 ;
      RECT 7.84 1.94 9.855 2.11 ;
      RECT 7.84 1.405 8.04 2.11 ;
      RECT 9.685 1.435 10.94 1.725 ;
      RECT 9.245 1.055 9.855 1.225 ;
      RECT 9.245 0.965 9.575 1.225 ;
      RECT 8.735 0.615 9.065 0.9 ;
      RECT 9.755 0.615 10.085 0.875 ;
      RECT 8.735 0.615 10.085 0.785 ;
      RECT 6.53 1.875 6.865 2.335 ;
      RECT 6.535 0.5 6.865 2.335 ;
      RECT 6.53 1.875 7.66 2.045 ;
      RECT 7.49 1.055 7.66 2.045 ;
      RECT 8.22 1.59 9.345 1.76 ;
      RECT 9.175 1.405 9.505 1.735 ;
      RECT 8.22 1.055 8.39 1.76 ;
      RECT 7.49 1.055 8.39 1.225 ;
      RECT 4.145 2.895 5.29 3.065 ;
      RECT 5.12 2.325 5.29 3.065 ;
      RECT 2.745 2.895 3.615 3.065 ;
      RECT 3.445 1.72 3.615 3.065 ;
      RECT 4.145 1.72 4.315 3.065 ;
      RECT 2.745 1.685 2.915 3.065 ;
      RECT 1.335 2 1.585 2.715 ;
      RECT 5.12 2.325 6.35 2.495 ;
      RECT 6.18 0.605 6.35 2.495 ;
      RECT 6.02 1.875 6.35 2.495 ;
      RECT 1.335 2 2.17 2.17 ;
      RECT 2 0.46 2.17 2.17 ;
      RECT 3.445 1.72 4.315 1.89 ;
      RECT 2 1.685 2.915 1.855 ;
      RECT 6.025 0.605 6.355 1.065 ;
      RECT 0.98 0.46 1.31 1.035 ;
      RECT 0.98 0.46 2.17 0.63 ;
      RECT 4.955 1.345 5.295 2.145 ;
      RECT 4.955 1.345 6 1.675 ;
      RECT 4.955 0.31 5.285 2.145 ;
      RECT 4.495 0.87 4.76 2.715 ;
      RECT 4.375 0.265 4.545 1.54 ;
      RECT 4.165 0.265 4.545 0.69 ;
      RECT 3.095 0.575 3.265 2.715 ;
      RECT 2.35 1.175 3.265 1.505 ;
      RECT 3.095 0.575 3.425 1.035 ;
      RECT 0.975 2.895 2.095 3.065 ;
      RECT 1.765 2.35 2.095 3.065 ;
      RECT 0.115 2.065 0.365 3.03 ;
      RECT 0.975 2.065 1.145 3.065 ;
      RECT 0.115 2.065 1.145 2.235 ;
  END
END scs130lp_sdfbbn_1

MACRO scs130lp_sdfbbn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfbbn_2 0 0 ;
  SIZE 18.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.87 1.11 4.2 1.78 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.495 0.81 1.795 1.795 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 17.365 0.265 17.695 3.065 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.485 1.815 15.765 3.065 ;
        RECT 15.595 0.265 15.765 3.065 ;
        RECT 15.41 0.265 15.765 1.125 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.525 1.345 14.92 1.78 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.215 0.55 1.885 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.895 1.215 1.315 1.885 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 0.932432 LAYER li ;
      ANTENNAMAXAREACAR 0.932432 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.851351 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.851351 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 12.575 1.18 12.865 1.41 ;
        RECT 8.255 1.225 12.865 1.365 ;
        RECT 8.255 1.18 8.545 1.41 ;
      LAYER li ;
        RECT 12.605 1.18 12.95 1.78 ;
        RECT 8.185 1.18 8.515 1.545 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 18.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 18.24 0.085 ;
        RECT 17.875 -0.085 18.125 1.095 ;
        RECT 16.935 -0.085 17.185 1.005 ;
        RECT 15.945 -0.085 16.195 1.125 ;
        RECT 14.98 -0.085 15.23 1.125 ;
        RECT 12.335 -0.085 12.665 0.65 ;
        RECT 10.205 -0.085 10.455 0.915 ;
        RECT 7.465 -0.085 7.795 0.65 ;
        RECT 5.38 -0.085 5.71 0.775 ;
        RECT 3.665 -0.085 3.995 0.915 ;
        RECT 2.325 -0.085 2.655 1.005 ;
        RECT 0.165 -0.085 0.495 1.035 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 18.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 18.24 3.415 ;
        RECT 17.875 1.815 18.125 3.415 ;
        RECT 16.935 1.815 17.185 3.415 ;
        RECT 15.945 1.815 16.195 3.415 ;
        RECT 14.975 2.74 15.305 3.415 ;
        RECT 13.935 2.74 14.265 3.415 ;
        RECT 12.685 2.47 12.935 3.415 ;
        RECT 9.51 1.875 9.84 3.415 ;
        RECT 7.955 2.425 8.285 3.415 ;
        RECT 5.36 2.675 5.69 3.415 ;
        RECT 3.645 2.385 3.895 3.415 ;
        RECT 2.72 2.425 3.05 3.415 ;
        RECT 0.77 2.415 1.1 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 16.425 0.295 16.755 2.64 ;
      RECT 16.425 1.185 17.185 1.515 ;
      RECT 13.115 2.12 13.445 3.065 ;
      RECT 13.115 2.39 15.305 2.56 ;
      RECT 15.135 1.305 15.305 2.56 ;
      RECT 13.665 0.995 13.835 2.56 ;
      RECT 12.23 2.12 13.445 2.29 ;
      RECT 12.23 1.96 12.56 2.29 ;
      RECT 15.135 1.305 15.415 1.635 ;
      RECT 13.48 0.615 13.81 1.165 ;
      RECT 14.015 1.96 14.795 2.21 ;
      RECT 14.015 0.995 14.34 2.21 ;
      RECT 14.015 0.995 14.8 1.165 ;
      RECT 14.47 0.665 14.8 1.165 ;
      RECT 13.99 0.265 14.24 0.815 ;
      RECT 12.925 0.265 13.255 0.65 ;
      RECT 12.925 0.265 14.24 0.435 ;
      RECT 11.03 2.12 11.47 2.715 ;
      RECT 11.3 0.575 11.47 2.715 ;
      RECT 13.13 1.46 13.485 1.79 ;
      RECT 13.13 0.83 13.3 1.79 ;
      RECT 11.3 0.575 11.63 1.255 ;
      RECT 11.3 0.83 13.3 1 ;
      RECT 10.68 2.895 12.02 3.065 ;
      RECT 11.69 1.7 12.02 3.065 ;
      RECT 10.68 1.095 10.85 3.065 ;
      RECT 10.68 1.095 11.12 1.675 ;
      RECT 6.77 0.83 6.945 1.545 ;
      RECT 9.855 1.095 11.12 1.265 ;
      RECT 9.855 0.265 10.025 1.265 ;
      RECT 6.77 0.83 8.145 1 ;
      RECT 7.975 0.265 8.145 1 ;
      RECT 7.975 0.265 10.025 0.435 ;
      RECT 8.525 2.075 9.33 2.755 ;
      RECT 9.16 1.055 9.33 2.755 ;
      RECT 7.475 2.075 9.33 2.245 ;
      RECT 7.475 1.825 7.655 2.245 ;
      RECT 10.17 1.445 10.5 1.705 ;
      RECT 9.16 1.445 10.5 1.615 ;
      RECT 8.835 0.965 9.165 1.225 ;
      RECT 8.325 0.615 8.655 1 ;
      RECT 9.345 0.615 9.675 0.875 ;
      RECT 8.325 0.615 9.675 0.785 ;
      RECT 6.42 2.075 6.75 2.755 ;
      RECT 6.42 2.075 7.295 2.245 ;
      RECT 7.125 1.475 7.295 2.245 ;
      RECT 6.42 0.665 6.59 2.755 ;
      RECT 7.835 1.725 8.98 1.895 ;
      RECT 8.705 1.405 8.98 1.895 ;
      RECT 7.835 1.475 8.005 1.895 ;
      RECT 7.125 1.475 8.005 1.645 ;
      RECT 4.075 2.895 5.18 3.065 ;
      RECT 5.01 2.325 5.18 3.065 ;
      RECT 4.075 2.035 4.245 3.065 ;
      RECT 5.91 2.295 6.24 2.755 ;
      RECT 6.07 0.665 6.24 2.755 ;
      RECT 1.65 2.035 1.98 2.715 ;
      RECT 5.01 2.325 6.24 2.495 ;
      RECT 1.65 2.035 4.245 2.205 ;
      RECT 1.975 0.46 2.145 2.205 ;
      RECT 5.91 0.665 6.24 1.125 ;
      RECT 0.985 0.46 1.315 1.035 ;
      RECT 0.985 0.46 2.145 0.63 ;
      RECT 4.95 0.315 5.2 2.145 ;
      RECT 4.95 1.815 5.89 1.985 ;
      RECT 5.615 1.315 5.89 1.985 ;
      RECT 4.87 0.315 5.2 0.775 ;
      RECT 4.425 1.005 4.77 2.715 ;
      RECT 4.425 0.455 4.595 2.715 ;
      RECT 4.175 0.455 4.595 0.915 ;
      RECT 2.325 1.515 3.445 1.855 ;
      RECT 2.945 0.575 3.445 1.855 ;
      RECT 2.325 1.185 2.58 1.855 ;
      RECT 1.3 2.895 2.49 3.065 ;
      RECT 2.16 2.385 2.49 3.065 ;
      RECT 0.26 2.065 0.59 3.065 ;
      RECT 1.3 2.065 1.47 3.065 ;
      RECT 0.26 2.065 1.47 2.235 ;
  END
END scs130lp_sdfbbn_2

MACRO scs130lp_sdfbbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfbbp_1 0 0 ;
  SIZE 15.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.445 1.5 3.775 2.17 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.465 1.525 1.795 1.855 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.38 1.815 15.75 3.065 ;
        RECT 15.58 0.265 15.75 3.065 ;
        RECT 15.38 0.265 15.75 1.125 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.96 1.765 14.315 3.065 ;
        RECT 14.145 0.265 14.315 3.065 ;
        RECT 13.88 0.265 14.315 1.075 ;
    END
  END QN
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.065 1.18 13.395 1.515 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.215 0.55 1.885 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.76 1.55 1.285 1.88 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 1.38536 LAYER li ;
      ANTENNAMAXAREACAR 1.38536 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.310811 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.310811 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 11.135 1.92 11.425 2.15 ;
        RECT 6.815 1.965 11.425 2.105 ;
        RECT 6.815 1.92 7.105 2.15 ;
      LAYER li ;
        RECT 11.08 1.765 11.41 2.15 ;
        RECT 6.995 1.375 7.525 1.78 ;
        RECT 6.845 1.95 7.165 2.15 ;
        RECT 6.995 1.375 7.165 2.15 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.84 0.085 ;
        RECT 14.95 -0.085 15.2 1.125 ;
        RECT 13.45 -0.085 13.7 1 ;
        RECT 10.86 -0.085 11.19 0.82 ;
        RECT 8.935 -0.085 9.265 0.595 ;
        RECT 7.005 -0.085 7.255 0.845 ;
        RECT 5.225 -0.085 5.475 0.65 ;
        RECT 3.265 -0.085 3.435 0.97 ;
        RECT 1.785 -0.085 2.035 0.995 ;
        RECT 0.175 -0.085 0.505 1.035 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.84 3.415 ;
        RECT 14.95 1.815 15.2 3.415 ;
        RECT 13.45 2.68 13.78 3.415 ;
        RECT 12.37 2.68 12.7 3.415 ;
        RECT 11.01 2.68 11.34 3.415 ;
        RECT 8.375 2.31 8.705 3.415 ;
        RECT 6.955 2.68 7.285 3.415 ;
        RECT 5.045 2.265 5.375 3.415 ;
        RECT 3.545 2.35 3.875 3.415 ;
        RECT 2.555 2.385 2.805 3.415 ;
        RECT 0.625 2.415 0.955 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 9.695 1.18 9.985 1.41 ;
      RECT 4.895 1.18 5.185 1.41 ;
      RECT 4.895 1.225 9.985 1.365 ;
    LAYER li ;
      RECT 14.52 0.665 14.77 2.495 ;
      RECT 14.52 1.305 15.4 1.635 ;
      RECT 11.52 2.33 11.85 3.065 ;
      RECT 10.575 2.33 13.78 2.5 ;
      RECT 13.61 1.255 13.78 2.5 ;
      RECT 12.15 1.205 12.32 2.5 ;
      RECT 10.575 1.745 10.87 2.5 ;
      RECT 13.61 1.255 13.965 1.585 ;
      RECT 11.94 1.205 12.32 1.535 ;
      RECT 12.94 1.765 13.27 2.15 ;
      RECT 12.5 1.765 13.27 1.935 ;
      RECT 12.5 0.83 12.8 1.935 ;
      RECT 8.525 0.775 8.82 1.315 ;
      RECT 10.485 1 11.76 1.17 ;
      RECT 13.02 0.635 13.27 1 ;
      RECT 11.59 0.83 13.27 1 ;
      RECT 10.485 0.265 10.655 1.17 ;
      RECT 8.525 0.775 9.615 0.945 ;
      RECT 9.445 0.265 9.615 0.945 ;
      RECT 9.445 0.265 10.655 0.435 ;
      RECT 12.4 0.265 12.65 0.65 ;
      RECT 11.37 0.265 11.7 0.65 ;
      RECT 11.37 0.265 12.65 0.435 ;
      RECT 9.28 2.595 9.61 3.015 ;
      RECT 9.28 2.595 10.395 2.765 ;
      RECT 10.225 1.35 10.395 2.765 ;
      RECT 11.59 1.715 11.97 2.045 ;
      RECT 11.59 1.35 11.76 2.045 ;
      RECT 10.135 1.35 11.76 1.52 ;
      RECT 10.135 0.615 10.305 1.52 ;
      RECT 9.795 0.615 10.305 0.945 ;
      RECT 9.61 2.085 10.045 2.415 ;
      RECT 9.61 1.125 9.955 2.415 ;
      RECT 7.465 1.96 7.795 2.725 ;
      RECT 6.485 2.33 7.795 2.5 ;
      RECT 6.485 1.45 6.655 2.5 ;
      RECT 7.465 1.96 9.36 2.13 ;
      RECT 9.03 1.125 9.36 2.13 ;
      RECT 8.175 0.645 8.345 2.13 ;
      RECT 6.485 1.45 6.815 1.77 ;
      RECT 7.945 0.645 8.345 0.815 ;
      RECT 7.435 0.265 7.765 0.845 ;
      RECT 7.435 0.265 8.705 0.465 ;
      RECT 6.135 0.265 6.305 2.725 ;
      RECT 7.705 1.025 7.995 1.695 ;
      RECT 6.135 1.025 7.995 1.195 ;
      RECT 6.135 0.265 6.465 1.195 ;
      RECT 5.625 2.265 5.955 2.725 ;
      RECT 5.785 0.265 5.955 2.725 ;
      RECT 1.485 2.035 1.815 2.715 ;
      RECT 1.485 2.035 2.145 2.205 ;
      RECT 1.975 1.175 2.145 2.205 ;
      RECT 0.995 1.175 2.385 1.345 ;
      RECT 2.215 0.265 2.385 1.345 ;
      RECT 2.915 1.15 3.785 1.32 ;
      RECT 3.615 0.265 3.785 1.32 ;
      RECT 0.995 0.575 1.325 1.345 ;
      RECT 2.915 0.265 3.085 1.32 ;
      RECT 4.875 0.83 5.955 1 ;
      RECT 5.705 0.265 5.955 1 ;
      RECT 4.875 0.265 5.045 1 ;
      RECT 3.615 0.265 5.045 0.435 ;
      RECT 2.215 0.265 3.085 0.435 ;
      RECT 4.525 1.915 4.865 2.945 ;
      RECT 4.525 1.915 5.56 2.085 ;
      RECT 5.045 1.415 5.56 2.085 ;
      RECT 4.525 0.615 4.695 2.945 ;
      RECT 5.045 1.18 5.215 2.085 ;
      RECT 4.925 1.18 5.215 1.41 ;
      RECT 4.055 0.615 4.345 3.03 ;
      RECT 3.965 0.615 4.345 1.73 ;
      RECT 2.985 2.385 3.315 3.065 ;
      RECT 2.985 1.685 3.155 3.065 ;
      RECT 2.325 1.685 3.155 1.855 ;
      RECT 2.325 1.525 2.735 1.855 ;
      RECT 2.565 0.615 2.735 1.855 ;
      RECT 1.135 2.895 2.325 3.065 ;
      RECT 1.995 2.385 2.325 3.065 ;
      RECT 0.115 2.065 0.445 3.065 ;
      RECT 1.135 2.065 1.305 3.065 ;
      RECT 0.115 2.065 1.305 2.235 ;
  END
END scs130lp_sdfbbp_1

MACRO scs130lp_sdfrbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrbp_1 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.41 1.2 4.645 1.78 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.475 0.78 1.805 1.525 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.475 0.355 12.82 2.285 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.4 1.855 13.765 3.075 ;
        RECT 13.585 0.355 13.765 3.075 ;
        RECT 13.395 0.355 13.765 1.175 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.555 1.155 2.86 2.215 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 1.695 2.385 1.865 ;
        RECT 2.07 1.395 2.385 1.865 ;
        RECT 0.555 1.535 1.305 1.865 ;
    END
  END SCE
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.411 LAYER met1 ;
      ANTENNAMAXAREACAR 1.479762 LAYER li ;
      ANTENNAMAXAREACAR 1.479762 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.420635 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.420635 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 10.175 1.92 10.465 2.15 ;
        RECT 3.455 1.965 10.465 2.105 ;
        RECT 7.775 1.92 8.065 2.15 ;
        RECT 3.455 1.92 3.745 2.15 ;
      LAYER li ;
        RECT 10.23 1.87 10.795 2.2 ;
        RECT 7.775 1.82 8.08 2.165 ;
        RECT 3.38 1.95 3.75 2.28 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.92 0.085 ;
        RECT 12.99 -0.085 13.225 1.175 ;
        RECT 11.545 -0.085 11.875 0.555 ;
        RECT 10.135 -0.085 10.465 0.61 ;
        RECT 7.95 -0.085 8.28 0.55 ;
        RECT 5.655 -0.085 5.835 0.96 ;
        RECT 4.665 -0.085 4.995 0.69 ;
        RECT 3.275 -0.085 3.605 0.655 ;
        RECT 0.585 -0.085 0.795 0.685 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.92 3.415 ;
        RECT 12.9 2.795 13.23 3.415 ;
        RECT 11.305 2.025 11.635 3.415 ;
        RECT 10.35 2.545 10.61 3.415 ;
        RECT 8.25 1.875 8.48 3.415 ;
        RECT 7.075 2.695 7.405 3.415 ;
        RECT 4.665 2.79 4.995 3.415 ;
        RECT 2.775 2.79 3.105 3.415 ;
        RECT 1.09 2.435 1.35 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 11.97 2.455 12.3 3.075 ;
      RECT 11.97 2.455 13.23 2.625 ;
      RECT 13.04 1.345 13.23 2.625 ;
      RECT 13.04 1.345 13.415 1.675 ;
      RECT 11.805 1.615 12.305 2.285 ;
      RECT 12.045 0.28 12.305 2.285 ;
      RECT 10.79 2.37 11.135 2.92 ;
      RECT 10.965 1.685 11.135 2.92 ;
      RECT 10.965 1.685 11.59 1.855 ;
      RECT 11.36 0.725 11.59 1.855 ;
      RECT 10 0.995 10.34 1.345 ;
      RECT 10 0.995 10.805 1.165 ;
      RECT 10.635 0.725 10.805 1.165 ;
      RECT 10.635 0.725 11.59 0.975 ;
      RECT 11.025 0.51 11.355 0.975 ;
      RECT 9.19 2.495 10.06 2.92 ;
      RECT 9.89 1.515 10.06 2.92 ;
      RECT 9.55 1.515 10.06 1.725 ;
      RECT 9.55 1.515 10.68 1.685 ;
      RECT 10.975 1.145 11.19 1.515 ;
      RECT 10.51 1.345 11.19 1.515 ;
      RECT 9.55 0.33 9.83 1.725 ;
      RECT 9.425 0.33 9.83 0.935 ;
      RECT 9.54 1.95 9.72 2.32 ;
      RECT 9.085 1.95 9.72 2.26 ;
      RECT 5.165 1.885 5.48 2.215 ;
      RECT 6.005 0.255 6.175 1.97 ;
      RECT 9.085 1.09 9.35 2.26 ;
      RECT 5.32 1.74 6.175 1.97 ;
      RECT 5.4 1.13 6.175 1.97 ;
      RECT 5.345 1.13 6.175 1.295 ;
      RECT 5.29 1.13 6.175 1.235 ;
      RECT 5.185 0.68 5.485 1.175 ;
      RECT 5.185 1.085 5.535 1.175 ;
      RECT 9.085 0.72 9.255 2.26 ;
      RECT 7.61 0.72 9.255 0.89 ;
      RECT 7.61 0.255 7.78 0.89 ;
      RECT 6.005 0.255 7.78 0.425 ;
      RECT 8.66 1.875 8.915 2.92 ;
      RECT 8.745 1.06 8.915 2.92 ;
      RECT 7.065 1.11 7.245 2.155 ;
      RECT 7.105 1.06 8.915 1.295 ;
      RECT 6.205 2.495 6.905 2.775 ;
      RECT 7.585 2.335 7.99 2.685 ;
      RECT 7.425 1.465 7.605 2.525 ;
      RECT 6.725 2.335 7.99 2.525 ;
      RECT 6.725 0.65 6.895 2.775 ;
      RECT 7.425 1.465 8.575 1.65 ;
      RECT 6.725 0.65 6.945 0.98 ;
      RECT 3.275 2.45 3.605 3.075 ;
      RECT 1.81 2.385 2.14 3.075 ;
      RECT 5.775 2.155 6.035 2.685 ;
      RECT 1.81 2.45 6.035 2.62 ;
      RECT 1.81 2.415 3.275 2.62 ;
      RECT 1.81 2.385 3.21 2.62 ;
      RECT 3.04 0.815 3.21 2.62 ;
      RECT 5.775 2.155 6.515 2.325 ;
      RECT 6.345 0.7 6.515 2.325 ;
      RECT 1.985 0.815 3.21 0.985 ;
      RECT 1.985 0.595 2.315 0.985 ;
      RECT 4.235 1.95 4.995 2.215 ;
      RECT 4.825 0.86 4.995 2.215 ;
      RECT 4.825 1.345 5.15 1.715 ;
      RECT 4.825 1.425 5.23 1.595 ;
      RECT 4.255 0.86 4.995 1.03 ;
      RECT 4.255 0.67 4.425 1.03 ;
      RECT 1.045 0.255 1.305 0.735 ;
      RECT 2.775 0.255 3.105 0.645 ;
      RECT 1.045 0.255 3.105 0.425 ;
      RECT 0.59 2.035 0.92 3.075 ;
      RECT 0.155 2.035 2.375 2.215 ;
      RECT 0.155 0.485 0.325 2.215 ;
      RECT 0.155 0.905 1.235 1.235 ;
      RECT 0.155 0.485 0.365 1.235 ;
  END
END scs130lp_sdfrbp_1

MACRO scs130lp_sdfrbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrbp_2 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.315 1.21 4.175 1.75 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.57 0.84 1.805 1.495 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.575 0.255 13.81 3.075 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.65 0.255 11.915 3.075 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.565 2.805 2.275 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.185 1.135 2.515 1.395 ;
        RECT 0.535 1.675 2.355 1.845 ;
        RECT 2.185 1.135 2.355 1.845 ;
        RECT 0.535 1.515 1.345 1.845 ;
    END
  END SCE
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.411 LAYER met1 ;
      ANTENNAMAXAREACAR 1.085714 LAYER li ;
      ANTENNAMAXAREACAR 1.085714 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.174603 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.174603 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 10.145 1.92 10.435 2.15 ;
        RECT 3.455 1.965 10.435 2.105 ;
        RECT 7.295 1.92 7.585 2.15 ;
        RECT 3.455 1.92 3.745 2.15 ;
      LAYER li ;
        RECT 10.125 1.94 10.505 2.3 ;
        RECT 7.3 1.825 7.605 2.155 ;
        RECT 3.325 1.92 3.695 2.2 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 14.4 0.085 ;
        RECT 13.98 -0.085 14.285 1.14 ;
        RECT 13.095 -0.085 13.405 1.06 ;
        RECT 12.085 -0.085 12.405 1.095 ;
        RECT 11.19 -0.085 11.48 0.9 ;
        RECT 9.88 -0.085 10.21 0.67 ;
        RECT 7.595 -0.085 7.925 0.55 ;
        RECT 5.26 -0.085 5.43 0.905 ;
        RECT 4.26 -0.085 4.59 0.69 ;
        RECT 3.35 -0.085 3.61 0.78 ;
        RECT 0.525 -0.085 0.855 0.765 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 14.4 3.415 ;
        RECT 13.98 1.815 14.285 3.415 ;
        RECT 13.095 1.815 13.405 3.415 ;
        RECT 12.085 1.795 12.405 3.415 ;
        RECT 11.15 2.28 11.48 3.415 ;
        RECT 9.71 2.85 10.455 3.415 ;
        RECT 10.105 2.525 10.455 3.415 ;
        RECT 7.775 2.085 8.025 3.415 ;
        RECT 6.69 2.675 7.02 3.415 ;
        RECT 4.215 2.825 4.545 3.415 ;
        RECT 2.67 2.835 3 3.415 ;
        RECT 1.05 2.435 1.31 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 12.575 0.285 12.885 2.495 ;
      RECT 12.575 1.23 13.405 1.56 ;
      RECT 12.575 0.285 12.905 1.56 ;
      RECT 10.625 2.47 10.895 2.855 ;
      RECT 10.675 1.94 10.895 2.855 ;
      RECT 10.675 1.94 11.235 2.11 ;
      RECT 11.065 1.07 11.235 2.11 ;
      RECT 10.125 1.07 11.235 1.26 ;
      RECT 9.615 0.86 11 1.19 ;
      RECT 10.67 0.33 11 1.26 ;
      RECT 8.825 2.49 9.155 2.91 ;
      RECT 8.825 2.49 9.935 2.67 ;
      RECT 9.765 1.36 9.935 2.67 ;
      RECT 8.825 2.08 9.105 2.91 ;
      RECT 9.765 1.43 10.875 1.76 ;
      RECT 9.24 1.36 9.955 1.53 ;
      RECT 9.24 0.255 9.445 1.53 ;
      RECT 9.02 0.255 9.445 0.65 ;
      RECT 9.275 1.99 9.595 2.32 ;
      RECT 4.685 1.815 5.085 2.315 ;
      RECT 4.95 1.05 5.12 2.145 ;
      RECT 9.275 1.7 9.515 2.32 ;
      RECT 8.73 1.7 9.515 1.9 ;
      RECT 4.95 1.075 5.77 1.78 ;
      RECT 5.6 0.31 5.77 1.78 ;
      RECT 8.73 0.82 9.07 1.9 ;
      RECT 4.905 1.075 5.77 1.155 ;
      RECT 4.77 0.595 5.09 1.11 ;
      RECT 8.705 0.82 9.07 0.965 ;
      RECT 8.67 0.82 9.07 0.93 ;
      RECT 7.245 0.72 8.85 0.89 ;
      RECT 7.245 0.775 8.9 0.89 ;
      RECT 7.245 0.31 7.425 0.89 ;
      RECT 5.6 0.31 7.425 0.48 ;
      RECT 8.31 2.08 8.63 2.91 ;
      RECT 6.62 1.06 6.79 2.155 ;
      RECT 8.31 1.06 8.56 2.91 ;
      RECT 6.62 1.06 8.56 1.235 ;
      RECT 7.19 2.335 7.565 2.695 ;
      RECT 5.795 2.335 6.52 2.695 ;
      RECT 5.795 2.335 7.565 2.505 ;
      RECT 6.96 1.405 7.13 2.505 ;
      RECT 5.795 2.29 6.45 2.695 ;
      RECT 6.28 0.65 6.45 2.695 ;
      RECT 7.965 1.405 8.14 1.735 ;
      RECT 6.96 1.405 8.14 1.645 ;
      RECT 6.28 0.65 6.62 0.89 ;
      RECT 3.21 2.485 3.54 3.075 ;
      RECT 1.77 2.445 2.1 3.075 ;
      RECT 1.77 2.485 5.625 2.655 ;
      RECT 5.39 1.95 5.625 2.655 ;
      RECT 5.355 2.325 5.625 2.655 ;
      RECT 1.77 2.445 3.145 2.655 ;
      RECT 2.975 0.795 3.145 2.655 ;
      RECT 5.39 1.95 6.11 2.12 ;
      RECT 5.94 0.65 6.11 2.12 ;
      RECT 1.975 0.795 3.145 0.965 ;
      RECT 1.975 0.605 2.305 0.965 ;
      RECT 3.865 1.93 4.115 2.315 ;
      RECT 3.865 1.93 4.515 2.1 ;
      RECT 4.345 0.86 4.515 2.1 ;
      RECT 4.345 1.28 4.78 1.61 ;
      RECT 3.8 0.86 4.515 1.04 ;
      RECT 3.8 0.595 4.06 1.04 ;
      RECT 1.115 0.265 1.415 0.765 ;
      RECT 1.115 0.265 1.49 0.685 ;
      RECT 2.85 0.265 3.18 0.625 ;
      RECT 1.115 0.265 3.18 0.435 ;
      RECT 0.53 2.015 0.88 3.075 ;
      RECT 0.53 2.015 2.335 2.265 ;
      RECT 0.095 2.015 2.335 2.195 ;
      RECT 0.095 0.935 0.365 2.195 ;
      RECT 0.095 0.935 1.255 1.265 ;
      RECT 0.095 0.465 0.355 2.195 ;
  END
END scs130lp_sdfrbp_2

MACRO scs130lp_sdfrbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrbp_lp 0 0 ;
  SIZE 19.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.43 1.295 15.76 1.78 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 0.265 3.235 0.67 ;
        RECT 1.78 0.265 3.235 0.435 ;
        RECT 1.78 0.265 2.11 0.535 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 18.755 0.265 19.085 3.065 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 16.5 1.765 16.83 3.065 ;
        RECT 16.66 0.265 16.83 3.065 ;
        RECT 16.445 0.265 16.83 1.075 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.335 1.55 3.685 1.965 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.477 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.475 1.18 0.805 2.15 ;
    END
  END SCE
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.189 LAYER li ;
      ANTENNAGATEAREA 0.633 LAYER met1 ;
      ANTENNAMAXAREACAR 1.355556 LAYER li ;
      ANTENNAMAXAREACAR 1.355556 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.089947 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.089947 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.15291 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 14.015 2.29 14.305 2.52 ;
        RECT 3.935 2.335 14.305 2.475 ;
        RECT 6.815 2.29 7.105 2.52 ;
        RECT 3.935 2.29 4.225 2.52 ;
      LAYER li ;
        RECT 13.665 2.1 14.275 2.52 ;
        RECT 6.755 2.225 7.085 2.52 ;
        RECT 3.865 1.625 4.195 2.52 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 19.2 0.245 ;
      LAYER li ;
        RECT 0 -0.085 19.2 0.085 ;
        RECT 17.965 -0.085 18.295 1.125 ;
        RECT 15.71 -0.085 16.04 0.71 ;
        RECT 12.18 -0.085 12.51 0.87 ;
        RECT 8.865 -0.085 9.195 0.465 ;
        RECT 6.995 -0.085 7.245 0.535 ;
        RECT 3.48 -0.085 3.65 0.555 ;
        RECT 0.945 -0.085 1.275 0.535 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 19.2 3.575 ;
      LAYER li ;
        RECT 0 3.245 19.2 3.415 ;
        RECT 17.965 1.815 18.295 3.415 ;
        RECT 15.71 1.96 16.04 3.415 ;
        RECT 13.93 2.7 14.18 3.415 ;
        RECT 12.495 2.795 12.825 3.415 ;
        RECT 8.895 1.855 9.225 3.415 ;
        RECT 5.86 2.735 6.19 3.415 ;
        RECT 2.895 2.495 3.225 3.415 ;
        RECT 0.96 2.495 1.29 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 17.06 0.665 17.39 2.495 ;
      RECT 17.06 1.305 18.575 1.635 ;
      RECT 10.93 2.425 11.26 2.715 ;
      RECT 10.93 2.425 11.96 2.595 ;
      RECT 11.79 0.575 11.96 2.595 ;
      RECT 11.79 1.745 13.05 1.915 ;
      RECT 12.72 1.4 13.05 1.915 ;
      RECT 16.015 1.255 16.345 1.585 ;
      RECT 12.72 1.4 14.49 1.57 ;
      RECT 14.32 0.89 14.49 1.57 ;
      RECT 14.055 1.24 14.49 1.57 ;
      RECT 16.015 0.89 16.185 1.585 ;
      RECT 14.32 0.89 16.185 1.06 ;
      RECT 11.13 0.575 11.96 0.905 ;
      RECT 14.5 0.265 15.25 0.71 ;
      RECT 12.69 0.265 13.02 0.595 ;
      RECT 12.69 0.265 15.25 0.435 ;
      RECT 14.92 1.24 15.25 3.065 ;
      RECT 14.685 1.24 15.25 1.57 ;
      RECT 14.36 2.7 14.69 3.03 ;
      RECT 14.52 1.75 14.69 3.03 ;
      RECT 12.595 2.095 13.4 2.265 ;
      RECT 13.23 1.75 13.4 2.265 ;
      RECT 13.23 1.75 14.69 1.92 ;
      RECT 12.14 1.05 12.47 1.565 ;
      RECT 12.14 1.05 12.86 1.22 ;
      RECT 13.89 0.685 14.14 1.06 ;
      RECT 12.69 0.89 14.14 1.06 ;
      RECT 13.14 2.445 13.47 3.03 ;
      RECT 12.14 2.445 13.47 2.615 ;
      RECT 12.14 2.185 12.415 2.615 ;
      RECT 10.465 2.895 12.315 3.065 ;
      RECT 11.985 2.795 12.315 3.065 ;
      RECT 10.465 2.295 10.715 3.065 ;
      RECT 9.415 2.895 10.285 3.065 ;
      RECT 10.115 1.945 10.285 3.065 ;
      RECT 9.415 0.995 9.585 3.065 ;
      RECT 7.99 0.615 8.24 2.715 ;
      RECT 11.36 1.915 11.61 2.245 ;
      RECT 10.115 1.945 11.61 2.115 ;
      RECT 11.08 1.915 11.61 2.115 ;
      RECT 11.08 1.085 11.25 2.115 ;
      RECT 6.185 1.065 6.515 1.375 ;
      RECT 10.62 1.085 11.25 1.255 ;
      RECT 6.185 1.065 8.24 1.235 ;
      RECT 7.85 0.615 8.24 1.235 ;
      RECT 7.85 0.995 9.585 1.165 ;
      RECT 10.62 0.575 10.95 1.255 ;
      RECT 9.765 0.265 9.935 2.715 ;
      RECT 9.765 1.435 10.9 1.765 ;
      RECT 9.765 0.265 10.095 1.765 ;
      RECT 6.57 0.715 7.67 0.885 ;
      RECT 7.5 0.265 7.67 0.885 ;
      RECT 8.42 0.645 10.095 0.815 ;
      RECT 4.38 0.265 4.71 0.715 ;
      RECT 6.57 0.265 6.74 0.885 ;
      RECT 8.42 0.265 8.59 0.815 ;
      RECT 7.5 0.265 8.59 0.435 ;
      RECT 4.38 0.265 6.74 0.435 ;
      RECT 7.64 2.895 8.59 3.065 ;
      RECT 8.42 1.345 8.59 3.065 ;
      RECT 7.64 1.885 7.81 3.065 ;
      RECT 5.855 1.885 6.155 2.215 ;
      RECT 5.855 1.885 7.81 2.055 ;
      RECT 8.42 1.345 9.235 1.675 ;
      RECT 7.21 2.7 7.46 3.065 ;
      RECT 4.715 2.385 4.905 2.895 ;
      RECT 6.37 2.7 7.46 2.87 ;
      RECT 6.37 2.385 6.54 2.87 ;
      RECT 4.715 2.385 6.54 2.555 ;
      RECT 5.505 1.235 5.675 2.555 ;
      RECT 5.505 1.545 7.81 1.715 ;
      RECT 7.48 1.415 7.81 1.715 ;
      RECT 4.53 1.235 4.86 1.535 ;
      RECT 4.53 1.235 5.675 1.405 ;
      RECT 4.1 1.075 4.35 1.445 ;
      RECT 4.18 0.885 4.35 1.445 ;
      RECT 4.18 0.885 5.77 1.055 ;
      RECT 5.47 0.715 6.39 0.885 ;
      RECT 2.075 2.145 2.405 3.065 ;
      RECT 3.405 2.7 4.545 2.975 ;
      RECT 4.375 2.025 4.545 2.975 ;
      RECT 3.405 2.145 3.575 2.975 ;
      RECT 0.985 2.145 3.575 2.315 ;
      RECT 4.375 2.025 5.325 2.195 ;
      RECT 5.075 1.585 5.325 2.195 ;
      RECT 0.985 1.065 1.155 2.315 ;
      RECT 1.685 1.065 2.015 1.615 ;
      RECT 0.985 1.065 2.015 1.235 ;
      RECT 2.475 1.065 2.725 1.615 ;
      RECT 2.475 1.065 3.585 1.235 ;
      RECT 3.415 0.725 3.585 1.235 ;
      RECT 3.415 0.725 4 0.895 ;
      RECT 3.83 0.265 4 0.895 ;
      RECT 3.83 0.265 4.21 0.715 ;
      RECT 1.335 1.795 3.155 1.965 ;
      RECT 2.905 1.415 3.155 1.965 ;
      RECT 1.335 1.415 1.505 1.965 ;
      RECT 0.125 2.435 0.5 3.065 ;
      RECT 0.125 0.265 0.295 3.065 ;
      RECT 0.125 0.715 2.68 0.885 ;
      RECT 2.295 0.615 2.68 0.885 ;
      RECT 0.125 0.265 0.455 0.885 ;
  END
END scs130lp_sdfrbp_lp

MACRO scs130lp_sdfrtn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrtn_1 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.475 1.345 4.645 1.75 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.51 1.07 2.885 1.405 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5817 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.88 1.815 13.345 3.075 ;
        RECT 13.085 0.295 13.345 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
      ANTENNAGATEAREA 0.411 LAYER met1 ;
      ANTENNAMAXAREACAR 6.372222 LAYER li ;
      ANTENNAMAXAREACAR 6.372222 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 5.472222 LAYER li ;
      ANTENNAMAXSIDEAREACAR 5.472222 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.181761 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.92 8.065 2.15 ;
        RECT 3.455 1.965 8.065 2.105 ;
        RECT 3.455 1.92 3.745 2.15 ;
      LAYER li ;
        RECT 10.145 1.375 11.04 1.965 ;
        RECT 9.095 2.905 10.315 3.075 ;
        RECT 10.145 1.375 10.315 3.075 ;
        RECT 9.095 2.635 9.265 3.075 ;
        RECT 8.545 2.635 9.265 2.805 ;
        RECT 8.545 1.43 8.715 2.805 ;
        RECT 7.755 1.43 8.715 1.745 ;
        RECT 7.755 1.43 8.025 2.18 ;
        RECT 3.46 1.525 3.695 2.195 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.64 0.745 1.885 1.955 ;
        RECT 0.95 0.745 1.885 1.095 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.055 1.575 2.785 1.85 ;
        RECT 2.055 1.575 2.62 2.105 ;
        RECT 2.055 1.055 2.34 2.105 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.44 0.085 ;
        RECT 12.525 -0.085 12.915 1.095 ;
        RECT 10.56 -0.085 10.89 0.855 ;
        RECT 8.12 -0.085 8.45 0.55 ;
        RECT 4.945 -0.085 5.275 0.455 ;
        RECT 3.875 -0.085 4.205 0.455 ;
        RECT 0.11 -0.085 0.405 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.44 3.415 ;
        RECT 12.37 2.585 12.71 3.415 ;
        RECT 12.45 1.765 12.71 3.415 ;
        RECT 11.55 2.71 11.84 3.415 ;
        RECT 10.54 2.71 10.87 3.415 ;
        RECT 8.585 2.985 8.915 3.415 ;
        RECT 7.155 2.69 7.455 3.415 ;
        RECT 4.945 2.77 5.275 3.415 ;
        RECT 3.755 2.77 4.085 3.415 ;
        RECT 1.955 2.955 2.625 3.415 ;
        RECT 0.11 1.815 0.405 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 11.81 2.135 12.28 2.415 ;
      RECT 12.11 0.35 12.28 2.415 ;
      RECT 12.11 1.265 12.915 1.595 ;
      RECT 12.11 0.35 12.355 1.595 ;
      RECT 11.08 2.175 11.38 3.075 ;
      RECT 10.495 2.175 11.39 2.505 ;
      RECT 11.22 1.795 11.39 2.505 ;
      RECT 11.22 1.795 11.94 1.965 ;
      RECT 11.77 0.595 11.94 1.965 ;
      RECT 11.465 0.595 11.94 0.855 ;
      RECT 9.63 2.405 9.965 2.735 ;
      RECT 9.795 0.625 9.965 2.735 ;
      RECT 11.34 1.025 11.6 1.495 ;
      RECT 9.62 0.625 9.965 1.295 ;
      RECT 9.62 1.025 11.6 1.205 ;
      RECT 5.395 1.815 6.16 2.26 ;
      RECT 5.395 1.815 6.63 2.15 ;
      RECT 9.28 1.755 9.625 2.085 ;
      RECT 5.395 0.965 5.82 2.26 ;
      RECT 9.28 0.255 9.45 2.085 ;
      RECT 5.395 1.125 6.63 1.295 ;
      RECT 6.46 0.255 6.63 1.295 ;
      RECT 7.18 0.72 9.45 0.89 ;
      RECT 9.195 0.255 9.45 0.89 ;
      RECT 7.18 0.255 7.35 0.89 ;
      RECT 6.46 0.255 7.35 0.51 ;
      RECT 9.195 0.255 10.11 0.455 ;
      RECT 8.94 2.265 9.46 2.465 ;
      RECT 8.94 1.06 9.11 2.465 ;
      RECT 7.215 1.06 7.545 2.145 ;
      RECT 7.215 1.06 9.11 1.26 ;
      RECT 7.625 2.35 8.375 3.02 ;
      RECT 8.195 1.985 8.375 3.02 ;
      RECT 6.405 2.32 6.695 3.02 ;
      RECT 6.405 2.35 8.375 2.52 ;
      RECT 6.405 2.32 7 2.52 ;
      RECT 6.8 0.68 7 2.52 ;
      RECT 3.195 2.365 3.525 3.065 ;
      RECT 5.915 2.43 6.235 3.02 ;
      RECT 1.105 2.615 1.435 2.965 ;
      RECT 1.105 2.615 3.525 2.785 ;
      RECT 3.195 2.43 6.235 2.6 ;
      RECT 3.195 2.365 4.035 2.6 ;
      RECT 3.865 0.625 4.035 2.6 ;
      RECT 6.04 0.625 6.29 0.955 ;
      RECT 2.255 0.685 4.035 0.855 ;
      RECT 3.865 0.625 6.29 0.795 ;
      RECT 2.255 0.605 2.585 0.855 ;
      RECT 4.32 1.93 5.215 2.26 ;
      RECT 5.045 0.965 5.215 2.26 ;
      RECT 4.385 0.965 5.215 1.165 ;
      RECT 1.35 0.265 1.68 0.545 ;
      RECT 3.22 0.265 3.55 0.515 ;
      RECT 1.35 0.265 3.55 0.435 ;
      RECT 0.575 1.815 0.81 2.495 ;
      RECT 0.575 2.275 2.96 2.445 ;
      RECT 2.79 2.02 2.96 2.445 ;
      RECT 0.575 1.965 1.425 2.445 ;
      RECT 2.79 2.02 3.265 2.195 ;
      RECT 3.095 1.035 3.265 2.195 ;
      RECT 0.575 0.295 0.77 2.495 ;
      RECT 3.095 1.035 3.425 1.205 ;
      RECT 0.575 0.295 0.87 0.565 ;
  END
END scs130lp_sdfrtn_1

MACRO scs130lp_sdfrtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrtp_1 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.55 1.425 11.88 2.5 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.565 2.255 1.805 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.085 0.255 13.355 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.411 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.94 2.255 9.27 2.57 ;
        RECT 8.035 2.475 9.215 2.645 ;
        RECT 6.77 2.905 8.285 3.075 ;
        RECT 8.035 2.475 8.285 3.075 ;
        RECT 6.77 2.32 6.95 3.075 ;
        RECT 5.8 2.32 6.95 2.49 ;
        RECT 5.8 1.94 6.13 2.545 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.965 1.175 3.31 2.145 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.54 1.2 2.795 1.395 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.44 0.085 ;
        RECT 12.575 -0.085 12.915 0.475 ;
        RECT 10.755 -0.085 11.085 0.475 ;
        RECT 8.49 -0.085 8.82 0.965 ;
        RECT 6.145 -0.085 6.475 0.615 ;
        RECT 3.405 -0.085 3.735 0.635 ;
        RECT 0.6 -0.085 0.895 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.44 3.415 ;
        RECT 12.43 2.015 12.915 3.415 ;
        RECT 10.715 2.71 11.04 3.415 ;
        RECT 9.79 2.71 10.05 3.415 ;
        RECT 8.455 2.855 9.19 3.415 ;
        RECT 6.27 2.66 6.6 3.415 ;
        RECT 4.865 2.505 5.195 3.415 ;
        RECT 3.04 2.655 3.37 3.415 ;
        RECT 1.32 2.315 1.65 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 10.175 1.18 10.465 1.41 ;
      RECT 7.295 1.18 7.585 1.41 ;
      RECT 4.895 1.18 5.185 1.41 ;
      RECT 3.935 1.18 4.225 1.41 ;
      RECT 3.935 1.225 10.465 1.365 ;
    LAYER li ;
      RECT 12.05 1.675 12.26 2.495 ;
      RECT 12.05 1.675 12.915 1.845 ;
      RECT 12.665 0.645 12.915 1.845 ;
      RECT 12.15 0.645 12.915 0.815 ;
      RECT 12.15 0.275 12.405 0.815 ;
      RECT 7.315 1.62 7.575 2.735 ;
      RECT 7.005 1.62 7.575 1.79 ;
      RECT 7.005 0.745 7.175 1.79 ;
      RECT 12.125 0.985 12.455 1.505 ;
      RECT 9.48 1.135 10.045 1.385 ;
      RECT 9.875 0.645 10.045 1.385 ;
      RECT 8.11 1.135 10.045 1.305 ;
      RECT 11.81 0.985 12.455 1.165 ;
      RECT 8.11 0.745 8.32 1.305 ;
      RECT 11.81 0.645 11.98 1.165 ;
      RECT 7.005 0.745 8.32 0.915 ;
      RECT 9.875 0.645 11.98 0.815 ;
      RECT 7.27 0.325 7.53 0.915 ;
      RECT 11.21 2.67 11.63 2.94 ;
      RECT 11.21 0.985 11.38 2.94 ;
      RECT 9.8 2.37 11.38 2.54 ;
      RECT 11.2 0.985 11.38 2.54 ;
      RECT 10.715 1.345 11.38 2.54 ;
      RECT 9.8 1.555 10.045 2.54 ;
      RECT 8.11 1.485 8.37 1.815 ;
      RECT 8.11 1.555 10.045 1.725 ;
      RECT 11.2 0.985 11.63 1.185 ;
      RECT 10.215 0.985 10.545 2.2 ;
      RECT 10.215 0.985 10.575 1.165 ;
      RECT 9.425 0.255 9.705 0.965 ;
      RECT 9.425 0.255 10.155 0.475 ;
      RECT 9.36 2.745 9.62 3.075 ;
      RECT 9.45 1.905 9.62 3.075 ;
      RECT 8.4 2.055 8.73 2.305 ;
      RECT 8.56 1.905 9.62 2.075 ;
      RECT 7.77 2.055 8.12 2.305 ;
      RECT 7.77 1.095 7.94 2.305 ;
      RECT 7.345 1.095 7.94 1.425 ;
      RECT 6.655 1.96 7.145 2.15 ;
      RECT 4.725 1.6 5.015 1.995 ;
      RECT 6.655 0.355 6.835 2.15 ;
      RECT 4.725 1.6 6.835 1.77 ;
      RECT 6.645 0.355 6.835 1.77 ;
      RECT 6.645 0.355 7.1 0.575 ;
      RECT 5.365 2.165 5.63 2.69 ;
      RECT 4.02 2.085 4.385 2.69 ;
      RECT 4.02 2.165 5.63 2.335 ;
      RECT 4.385 0.785 4.555 2.335 ;
      RECT 6.145 0.785 6.475 1.43 ;
      RECT 4.385 0.785 6.475 0.995 ;
      RECT 2.11 2.315 2.44 2.995 ;
      RECT 3.54 2.295 3.825 2.965 ;
      RECT 2.11 2.315 3.825 2.485 ;
      RECT 3.48 0.815 3.685 2.485 ;
      RECT 1.99 0.815 4.215 0.985 ;
      RECT 4.015 0.655 4.215 0.985 ;
      RECT 1.99 0.615 2.32 0.985 ;
      RECT 2.895 0.265 3.225 0.635 ;
      RECT 1.145 0.265 1.355 0.595 ;
      RECT 1.145 0.265 3.225 0.435 ;
      RECT 0.09 1.975 1.15 2.965 ;
      RECT 0.09 1.975 2.675 2.145 ;
      RECT 2.425 1.815 2.675 2.145 ;
      RECT 0.09 0.415 0.37 2.965 ;
      RECT 0.09 0.86 1.51 1.03 ;
      RECT 0.09 0.415 0.43 1.03 ;
      RECT 4.735 1.165 5.125 1.43 ;
      RECT 3.855 1.155 4.215 1.915 ;
  END
END scs130lp_sdfrtp_1

MACRO scs130lp_sdfrtp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrtp_2 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.63 1.415 12.005 2.49 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 1.55 2.735 1.76 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.115 1.755 13.375 3.075 ;
        RECT 13.2 0.255 13.375 3.075 ;
        RECT 13.115 0.255 13.375 1.065 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.411 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.755 2.525 9.405 2.695 ;
        RECT 9.075 2.25 9.405 2.695 ;
        RECT 6.755 2.305 6.925 2.695 ;
        RECT 5.795 2.305 6.925 2.475 ;
        RECT 5.795 1.95 6.125 2.475 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.905 1.21 3.285 2.13 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 1.2 2.735 1.38 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.92 0.085 ;
        RECT 13.545 -0.085 13.815 1.095 ;
        RECT 12.615 -0.085 12.945 0.475 ;
        RECT 10.88 -0.085 11.21 0.475 ;
        RECT 8.47 -0.085 8.8 0.955 ;
        RECT 6.145 -0.085 6.475 0.615 ;
        RECT 3.405 -0.085 3.735 0.665 ;
        RECT 0.565 -0.085 0.895 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.92 3.415 ;
        RECT 13.545 1.815 13.815 3.415 ;
        RECT 12.545 2.015 12.945 3.415 ;
        RECT 10.805 2.665 11.12 3.415 ;
        RECT 9.925 2.705 10.175 3.415 ;
        RECT 8.41 2.865 9.14 3.415 ;
        RECT 6.245 2.645 6.575 3.415 ;
        RECT 4.855 2.515 5.185 3.415 ;
        RECT 2.97 2.64 3.3 3.415 ;
        RECT 1.205 2.32 1.475 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 10.175 1.18 10.465 1.41 ;
      RECT 7.295 1.18 7.585 1.41 ;
      RECT 4.895 1.18 5.185 1.41 ;
      RECT 3.935 1.18 4.225 1.41 ;
      RECT 3.935 1.225 10.465 1.365 ;
    LAYER li ;
      RECT 12.175 1.675 12.375 2.495 ;
      RECT 12.175 1.675 12.89 1.845 ;
      RECT 12.72 0.645 12.89 1.845 ;
      RECT 12.72 1.245 13.03 1.575 ;
      RECT 12.72 0.645 12.945 1.575 ;
      RECT 12.275 0.645 12.945 0.815 ;
      RECT 12.275 0.275 12.445 0.815 ;
      RECT 12.115 0.275 12.445 0.465 ;
      RECT 7.27 1.605 7.555 2.355 ;
      RECT 7.005 1.605 7.555 1.775 ;
      RECT 7.005 0.325 7.175 1.775 ;
      RECT 12.21 0.995 12.54 1.505 ;
      RECT 8.065 1.205 10 1.375 ;
      RECT 9.83 0.645 10 1.375 ;
      RECT 11.9 0.995 12.54 1.245 ;
      RECT 8.065 0.325 8.235 1.375 ;
      RECT 11.9 0.645 12.07 1.245 ;
      RECT 7.005 0.325 8.235 0.925 ;
      RECT 9.83 0.645 12.07 0.815 ;
      RECT 11.29 2.66 11.72 2.94 ;
      RECT 11.29 0.985 11.46 2.94 ;
      RECT 9.935 2.325 11.46 2.495 ;
      RECT 10.805 1.345 11.46 2.495 ;
      RECT 9.935 1.56 10.105 2.495 ;
      RECT 8.065 1.56 8.325 1.885 ;
      RECT 8.065 1.56 10.105 1.73 ;
      RECT 8.065 1.555 8.245 1.885 ;
      RECT 11.29 0.985 11.72 1.245 ;
      RECT 10.375 0.985 10.635 2.155 ;
      RECT 10.21 0.985 10.635 1.425 ;
      RECT 10.21 0.985 10.7 1.165 ;
      RECT 9.38 0.255 9.66 0.97 ;
      RECT 9.38 0.255 10.11 0.475 ;
      RECT 9.31 2.865 9.755 3.075 ;
      RECT 9.585 1.91 9.755 3.075 ;
      RECT 8.535 1.91 8.865 2.275 ;
      RECT 8.535 1.91 9.755 2.08 ;
      RECT 7.725 2.095 8.075 2.355 ;
      RECT 7.725 1.095 7.895 2.355 ;
      RECT 7.345 1.095 7.895 1.425 ;
      RECT 6.655 1.945 7.1 2.135 ;
      RECT 4.725 1.6 5.01 1.995 ;
      RECT 6.655 0.325 6.835 2.135 ;
      RECT 4.725 1.6 6.835 1.77 ;
      RECT 6.645 0.325 6.835 1.77 ;
      RECT 5.355 2.175 5.625 2.695 ;
      RECT 4.055 2.175 4.385 2.695 ;
      RECT 4.055 2.175 5.625 2.345 ;
      RECT 4.385 0.64 4.555 2.345 ;
      RECT 6.145 0.785 6.475 1.43 ;
      RECT 4.385 0.785 6.475 0.995 ;
      RECT 4.385 0.64 4.8 0.995 ;
      RECT 1.995 2.3 2.325 3 ;
      RECT 3.51 2.3 3.885 2.97 ;
      RECT 1.995 2.3 3.885 2.47 ;
      RECT 3.455 0.835 3.68 2.47 ;
      RECT 1.99 0.835 4.215 1.005 ;
      RECT 3.955 0.64 4.215 1.005 ;
      RECT 1.99 0.605 2.32 1.005 ;
      RECT 2.895 0.265 3.225 0.665 ;
      RECT 1.085 0.265 1.415 0.625 ;
      RECT 1.085 0.265 3.225 0.435 ;
      RECT 0.135 1.93 1.035 3 ;
      RECT 0.135 1.93 2.56 2.13 ;
      RECT 0.135 0.86 0.405 3 ;
      RECT 0.135 0.86 1.51 1.03 ;
      RECT 0.135 0.415 0.395 3 ;
      RECT 4.735 1.165 5.2 1.43 ;
      RECT 3.85 1.175 4.215 1.995 ;
  END
END scs130lp_sdfrtp_2

MACRO scs130lp_sdfrtp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrtp_4 0 0 ;
  SIZE 15.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.155 1.525 12.57 2.525 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.05 1.57 2.325 1.76 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2096 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.665 1.735 15.26 1.985 ;
        RECT 15 1.055 15.26 1.985 ;
        RECT 13.665 1.055 15.26 1.225 ;
        RECT 13.665 1.045 14.79 1.225 ;
        RECT 14.525 0.255 14.79 1.225 ;
        RECT 14.545 1.735 14.745 3.075 ;
        RECT 13.665 1.735 13.875 3.075 ;
        RECT 13.665 0.255 13.855 1.225 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.411 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.19 2.485 9.69 2.655 ;
        RECT 9.36 2.245 9.69 2.655 ;
        RECT 7.2 2.725 8.36 2.895 ;
        RECT 8.19 2.485 8.36 2.895 ;
        RECT 7.2 2.285 7.37 2.895 ;
        RECT 6.41 2.285 7.37 2.455 ;
        RECT 6.41 1.895 6.58 2.455 ;
        RECT 6.21 1.895 6.58 2.13 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.025 1.29 3.475 2.125 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.55 1.205 2.805 1.4 ;
        RECT 0.55 1.205 0.88 1.76 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.36 0.085 ;
        RECT 14.96 -0.085 15.255 0.885 ;
        RECT 14.025 -0.085 14.355 0.875 ;
        RECT 13.165 -0.085 13.495 0.665 ;
        RECT 11.175 -0.085 11.505 0.455 ;
        RECT 8.955 -0.085 9.285 0.965 ;
        RECT 6.435 -0.085 6.765 0.995 ;
        RECT 3.355 -0.085 3.615 0.725 ;
        RECT 0.525 -0.085 0.855 0.625 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.36 3.415 ;
        RECT 14.925 2.155 15.255 3.415 ;
        RECT 14.045 2.155 14.375 3.415 ;
        RECT 13.165 2.095 13.495 3.415 ;
        RECT 11.095 2.665 11.61 3.415 ;
        RECT 11.43 2.105 11.61 3.415 ;
        RECT 10.21 2.665 10.41 3.415 ;
        RECT 9.005 2.825 9.335 3.415 ;
        RECT 6.69 2.625 7.02 3.415 ;
        RECT 5.36 2.475 5.7 3.415 ;
        RECT 3.355 2.645 3.685 3.415 ;
        RECT 1.62 2.295 1.91 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 10.655 1.18 10.945 1.41 ;
      RECT 7.775 1.18 8.065 1.41 ;
      RECT 5.375 1.18 5.665 1.41 ;
      RECT 4.415 1.18 4.705 1.41 ;
      RECT 4.415 1.225 10.945 1.365 ;
    LAYER li ;
      RECT 12.74 1.755 12.995 3.075 ;
      RECT 12.74 1.755 13.475 1.925 ;
      RECT 13.305 0.835 13.475 1.925 ;
      RECT 13.305 1.395 14.82 1.565 ;
      RECT 12.735 0.835 13.475 1.015 ;
      RECT 12.735 0.255 12.995 1.015 ;
      RECT 7.735 1.56 8.02 2.545 ;
      RECT 7.485 1.56 8.02 1.73 ;
      RECT 7.485 0.395 7.655 1.73 ;
      RECT 12.86 1.185 13.135 1.515 ;
      RECT 9.72 1.135 10.485 1.375 ;
      RECT 10.315 0.625 10.485 1.375 ;
      RECT 12.3 1.185 13.135 1.355 ;
      RECT 8.54 1.135 10.485 1.305 ;
      RECT 12.3 0.625 12.47 1.355 ;
      RECT 8.54 0.395 8.71 1.305 ;
      RECT 7.485 0.395 8.71 0.945 ;
      RECT 10.315 0.625 12.47 0.795 ;
      RECT 11.805 2.67 12.06 3 ;
      RECT 11.805 0.975 11.985 3 ;
      RECT 10.22 2.325 11.26 2.495 ;
      RECT 11.09 1.345 11.26 2.495 ;
      RECT 10.22 1.555 10.39 2.495 ;
      RECT 8.53 1.485 8.79 1.815 ;
      RECT 8.53 1.555 10.39 1.725 ;
      RECT 11.09 1.345 11.985 1.675 ;
      RECT 11.79 0.975 11.985 1.675 ;
      RECT 11.79 0.975 12.12 1.165 ;
      RECT 10.665 0.965 10.92 2.145 ;
      RECT 10.665 0.965 10.995 1.165 ;
      RECT 9.845 0.255 10.145 0.965 ;
      RECT 9.845 0.255 10.575 0.455 ;
      RECT 9.595 2.825 10.04 3.045 ;
      RECT 9.87 1.905 10.04 3.045 ;
      RECT 8.82 2.055 9.15 2.315 ;
      RECT 8.98 1.905 10.04 2.075 ;
      RECT 8.19 2.055 8.54 2.315 ;
      RECT 8.19 1.175 8.36 2.315 ;
      RECT 7.835 1.175 8.36 1.38 ;
      RECT 7.115 1.9 7.565 2.115 ;
      RECT 5.265 1.665 6.04 1.965 ;
      RECT 7.115 0.335 7.315 2.115 ;
      RECT 7.105 0.335 7.315 1.725 ;
      RECT 5.87 1.555 7.315 1.725 ;
      RECT 4.405 2.135 4.825 2.775 ;
      RECT 5.87 2.36 6.24 2.69 ;
      RECT 5.87 2.135 6.04 2.69 ;
      RECT 4.405 2.135 6.04 2.305 ;
      RECT 4.815 1.21 4.995 2.305 ;
      RECT 5.785 1.165 6.935 1.385 ;
      RECT 4.815 1.21 5.215 1.38 ;
      RECT 5.045 0.64 5.215 1.38 ;
      RECT 5.785 0.64 5.955 1.385 ;
      RECT 5.045 0.64 5.955 0.955 ;
      RECT 2.37 2.295 2.7 2.975 ;
      RECT 3.855 0.64 4.235 2.905 ;
      RECT 2.37 2.295 4.235 2.475 ;
      RECT 3.78 0.895 4.235 2.475 ;
      RECT 2.905 0.895 4.235 1.065 ;
      RECT 1.95 0.815 3.075 0.985 ;
      RECT 3.785 0.64 4.875 0.97 ;
      RECT 1.95 0.595 2.28 0.985 ;
      RECT 2.855 0.255 3.185 0.645 ;
      RECT 1.045 0.255 1.375 0.625 ;
      RECT 1.045 0.255 3.185 0.425 ;
      RECT 1.15 1.93 1.45 2.975 ;
      RECT 0.155 1.93 1.45 2.275 ;
      RECT 0.155 1.93 2.855 2.125 ;
      RECT 2.605 1.77 2.855 2.125 ;
      RECT 0.155 0.795 0.38 2.275 ;
      RECT 0.155 0.795 1.5 1.03 ;
      RECT 0.155 0.415 0.355 2.275 ;
      RECT 5.385 1.125 5.615 1.455 ;
      RECT 4.405 1.14 4.645 1.88 ;
  END
END scs130lp_sdfrtp_4

MACRO scs130lp_sdfrtp_lp2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrtp_lp2 0 0 ;
  SIZE 16.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.825 1.17 5.155 1.5 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.575 1.51 0.905 1.84 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.645 1.92 16.205 2.96 ;
        RECT 15.875 0.43 16.205 2.96 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.895 1.45 2.255 1.78 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 1.555 3.875 1.885 ;
        RECT 1.085 1.96 3.655 2.13 ;
        RECT 3.485 1.555 3.655 2.13 ;
        RECT 1.085 1.55 1.685 2.13 ;
    END
  END SCE
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
      ANTENNAGATEAREA 0.939 LAYER met1 ;
      ANTENNAMAXAREACAR 1.396645 LAYER li ;
      ANTENNAMAXAREACAR 1.396645 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.399361 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.399361 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.092332 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 12.575 1.55 12.865 1.78 ;
        RECT 2.975 1.595 12.865 1.735 ;
        RECT 8.735 1.55 9.025 1.78 ;
        RECT 2.975 1.55 3.265 1.78 ;
      LAYER li ;
        RECT 13.085 1.615 13.485 1.935 ;
        RECT 13.085 1.615 13.315 2.89 ;
        RECT 12.635 1.615 13.485 1.785 ;
        RECT 12.635 1.55 12.835 1.785 ;
        RECT 8.765 1.325 9.2 1.645 ;
        RECT 8.765 1.325 9.185 1.78 ;
        RECT 2.975 1.45 3.305 1.78 ;
    END
  END RESETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 16.32 0.085 ;
        RECT 15.085 -0.085 15.415 0.89 ;
        RECT 12.635 -0.085 12.965 0.51 ;
        RECT 8.85 -0.085 9.18 0.445 ;
        RECT 5.21 -0.085 5.54 0.725 ;
        RECT 2.56 -0.085 2.89 0.88 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 16.32 3.415 ;
        RECT 15.115 1.92 15.445 3.415 ;
        RECT 14.025 2.075 14.355 3.415 ;
        RECT 12.4 2.075 12.65 3.415 ;
        RECT 10.08 1.685 10.41 3.415 ;
        RECT 8.585 2.31 8.915 3.415 ;
        RECT 5.18 2.81 5.51 3.415 ;
        RECT 3.22 2.855 3.55 3.415 ;
        RECT 1.58 2.66 1.91 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 14.535 1.57 14.915 2.96 ;
      RECT 14.535 1.57 15.68 1.74 ;
      RECT 15.35 1.07 15.68 1.74 ;
      RECT 14.535 0.43 14.705 2.96 ;
      RECT 14.375 0.43 14.705 0.89 ;
      RECT 13.495 2.115 13.835 3.065 ;
      RECT 13.665 1.265 13.835 3.065 ;
      RECT 13.015 1.265 14.195 1.435 ;
      RECT 14.025 0.295 14.195 1.435 ;
      RECT 12.635 1.04 13.185 1.37 ;
      RECT 13.67 0.295 14.195 0.51 ;
      RECT 11.3 1.685 11.63 3.065 ;
      RECT 11.3 1.685 12.455 1.855 ;
      RECT 12.285 0.505 12.455 1.855 ;
      RECT 13.515 0.69 13.845 1.085 ;
      RECT 12.285 0.69 13.845 0.86 ;
      RECT 11.51 0.505 12.455 0.675 ;
      RECT 11.51 0.265 11.84 0.675 ;
      RECT 10.955 1.12 12.105 1.45 ;
      RECT 11.815 0.91 12.105 1.45 ;
      RECT 10.605 1.685 11.02 2.725 ;
      RECT 10.605 0.275 10.775 2.725 ;
      RECT 8.225 0.975 8.555 1.525 ;
      RECT 9.87 1.275 10.775 1.445 ;
      RECT 9.87 0.975 10.04 1.445 ;
      RECT 8.225 0.975 10.04 1.145 ;
      RECT 10.005 0.275 10.775 0.445 ;
      RECT 7.555 0.625 7.725 1.525 ;
      RECT 10.21 0.625 10.425 1.095 ;
      RECT 7.555 0.625 10.425 0.795 ;
      RECT 9.275 1.96 9.7 2.755 ;
      RECT 9.37 1.325 9.7 2.755 ;
      RECT 7.215 1.79 7.79 2.755 ;
      RECT 7.215 1.96 9.7 2.13 ;
      RECT 9.355 1.715 9.7 2.755 ;
      RECT 7.215 0.625 7.385 2.755 ;
      RECT 3.73 2.895 5.01 3.065 ;
      RECT 4.84 2.46 5.01 3.065 ;
      RECT 2.69 2.31 3.02 3.065 ;
      RECT 0.09 2.075 0.89 3.065 ;
      RECT 3.73 2.505 3.9 3.065 ;
      RECT 6.865 0.595 7.035 2.755 ;
      RECT 2.69 2.505 3.9 2.675 ;
      RECT 4.84 2.46 7.035 2.63 ;
      RECT 0.09 2.31 3.02 2.48 ;
      RECT 0.09 0.62 0.26 3.065 ;
      RECT 6.705 0.595 7.035 1.145 ;
      RECT 1.15 0.615 1.48 0.865 ;
      RECT 0.09 0.62 1.48 0.79 ;
      RECT 5.71 2.03 6.29 2.28 ;
      RECT 5.975 1.45 6.29 2.28 ;
      RECT 5.975 1.45 6.685 1.78 ;
      RECT 6.07 0.595 6.455 1.78 ;
      RECT 4.42 1.68 4.67 2.715 ;
      RECT 4.42 1.68 5.805 1.85 ;
      RECT 5.475 1.18 5.805 1.85 ;
      RECT 4.42 0.635 4.59 2.715 ;
      RECT 3.835 2.075 4.225 2.325 ;
      RECT 4.055 0.595 4.225 2.325 ;
      RECT 2.435 1.1 2.765 1.78 ;
      RECT 0.44 0.97 0.735 1.3 ;
      RECT 0.44 1.1 4.225 1.27 ;
      RECT 3.82 0.595 4.225 1.27 ;
      RECT 2.05 0.265 2.38 0.88 ;
      RECT 0.17 0.265 0.5 0.44 ;
      RECT 0.17 0.265 2.38 0.435 ;
  END
END scs130lp_sdfrtp_lp2

MACRO scs130lp_sdfrtp_ov2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfrtp_ov2 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.55 1.425 11.88 2.5 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.565 2.255 1.805 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.085 0.255 13.355 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.378 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.94 2.255 9.27 2.57 ;
        RECT 8.035 2.475 9.215 2.645 ;
        RECT 6.77 2.905 8.285 3.075 ;
        RECT 8.035 2.475 8.285 3.075 ;
        RECT 6.77 2.32 6.95 3.075 ;
        RECT 5.8 2.32 6.95 2.49 ;
        RECT 5.8 1.94 6.13 2.545 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.965 1.175 3.31 2.145 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.54 1.2 2.795 1.395 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.44 0.085 ;
        RECT 12.575 -0.085 12.915 0.475 ;
        RECT 10.755 -0.085 11.085 0.475 ;
        RECT 8.49 -0.085 8.82 0.965 ;
        RECT 6.145 -0.085 6.475 0.94 ;
        RECT 3.405 -0.085 3.735 0.635 ;
        RECT 0.6 -0.085 0.895 0.69 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.44 3.415 ;
        RECT 12.43 2.015 12.915 3.415 ;
        RECT 10.755 2.71 11.04 3.415 ;
        RECT 9.79 2.71 10.05 3.415 ;
        RECT 8.455 2.855 9.19 3.415 ;
        RECT 6.27 2.66 6.6 3.415 ;
        RECT 4.865 2.505 5.195 3.415 ;
        RECT 3.07 2.655 3.4 3.415 ;
        RECT 1.32 2.39 1.65 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 10.175 1.18 10.465 1.41 ;
      RECT 7.295 1.18 7.585 1.41 ;
      RECT 4.895 1.18 5.185 1.41 ;
      RECT 3.935 1.18 4.225 1.41 ;
      RECT 3.935 1.225 10.465 1.365 ;
    LAYER li ;
      RECT 12.05 1.675 12.26 2.495 ;
      RECT 12.05 1.675 12.915 1.845 ;
      RECT 12.665 0.645 12.915 1.845 ;
      RECT 12.15 0.645 12.915 0.815 ;
      RECT 12.15 0.275 12.405 0.815 ;
      RECT 7.315 1.62 7.575 2.735 ;
      RECT 7.005 1.62 7.575 1.79 ;
      RECT 7.005 0.745 7.175 1.79 ;
      RECT 12.125 0.985 12.455 1.505 ;
      RECT 9.48 1.135 10.045 1.385 ;
      RECT 9.875 0.645 10.045 1.385 ;
      RECT 8.11 1.135 10.045 1.305 ;
      RECT 11.81 0.985 12.455 1.165 ;
      RECT 8.11 0.745 8.32 1.305 ;
      RECT 11.81 0.645 11.98 1.165 ;
      RECT 7.005 0.745 8.32 0.915 ;
      RECT 9.875 0.645 11.98 0.815 ;
      RECT 7.2 0.625 7.87 0.915 ;
      RECT 11.21 2.715 11.63 3.045 ;
      RECT 11.21 0.985 11.38 3.045 ;
      RECT 9.8 2.37 11.38 2.54 ;
      RECT 11.2 0.985 11.38 2.54 ;
      RECT 10.715 1.345 11.38 2.54 ;
      RECT 9.8 1.555 10.045 2.54 ;
      RECT 8.11 1.485 8.37 1.815 ;
      RECT 8.11 1.555 10.045 1.725 ;
      RECT 11.2 0.985 11.63 1.185 ;
      RECT 10.215 0.985 10.545 2.2 ;
      RECT 10.215 0.985 10.575 1.165 ;
      RECT 9.425 0.255 9.705 0.965 ;
      RECT 9.425 0.255 10.155 0.475 ;
      RECT 9.36 2.745 9.62 3.075 ;
      RECT 9.45 1.905 9.62 3.075 ;
      RECT 8.4 2.055 8.73 2.305 ;
      RECT 8.56 1.905 9.62 2.075 ;
      RECT 7.77 2.055 8.12 2.305 ;
      RECT 7.77 1.095 7.94 2.305 ;
      RECT 7.345 1.095 7.94 1.425 ;
      RECT 6.655 1.96 7.145 2.15 ;
      RECT 4.725 1.6 5.015 1.995 ;
      RECT 6.655 0.63 6.835 2.15 ;
      RECT 4.725 1.6 6.835 1.77 ;
      RECT 6.645 0.63 6.835 1.77 ;
      RECT 5.365 2.165 5.63 2.69 ;
      RECT 4.065 2.085 4.385 2.69 ;
      RECT 4.065 2.165 5.63 2.335 ;
      RECT 4.385 0.785 4.555 2.335 ;
      RECT 5.465 1.17 6.475 1.43 ;
      RECT 5.465 0.785 5.67 1.43 ;
      RECT 4.385 0.785 5.67 0.995 ;
      RECT 2.11 2.315 2.44 2.68 ;
      RECT 3.59 2.295 3.885 2.625 ;
      RECT 2.11 2.315 3.885 2.485 ;
      RECT 3.48 0.815 3.685 2.485 ;
      RECT 1.99 0.815 4.215 0.985 ;
      RECT 4.015 0.655 4.215 0.985 ;
      RECT 1.99 0.615 2.32 0.985 ;
      RECT 2.895 0.265 3.225 0.635 ;
      RECT 1.145 0.265 1.355 0.595 ;
      RECT 1.145 0.265 3.225 0.435 ;
      RECT 0.09 1.975 1.14 2.965 ;
      RECT 0.09 1.975 2.675 2.145 ;
      RECT 2.425 1.815 2.675 2.145 ;
      RECT 0.09 0.415 0.37 2.965 ;
      RECT 0.09 0.86 1.51 1.03 ;
      RECT 0.09 0.415 0.43 1.03 ;
      RECT 4.735 1.165 5.125 1.43 ;
      RECT 3.855 1.155 4.215 1.915 ;
  END
END scs130lp_sdfrtp_ov2

MACRO scs130lp_sdfsbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfsbp_1 0 0 ;
  SIZE 15.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.275 0.83 3.755 1.885 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.105 0.765 1.915 1.775 ;
        RECT 1.105 0.765 1.555 1.945 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5733 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.915 1.02 14.25 3.075 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.835 1.84 15.275 3.075 ;
        RECT 15.005 0.38 15.275 3.075 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.08 2.735 2.205 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.56 2.125 2.375 2.295 ;
        RECT 2.125 0.995 2.375 2.295 ;
        RECT 0.56 1.915 0.935 2.295 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.252 LAYER met1 ;
      ANTENNAMAXAREACAR 1.466667 LAYER li ;
      ANTENNAMAXAREACAR 1.466667 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.730159 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.730159 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 10.655 1.92 10.945 2.15 ;
        RECT 7.295 1.965 10.945 2.105 ;
        RECT 7.295 1.92 7.585 2.15 ;
      LAYER li ;
        RECT 10.65 1.92 11.53 2.13 ;
        RECT 7.345 1.79 7.645 2.13 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.36 0.085 ;
        RECT 14.425 -0.085 14.755 0.51 ;
        RECT 11.9 -0.085 12.455 1.08 ;
        RECT 10.82 -0.085 11.15 0.96 ;
        RECT 8.855 -0.085 9.055 0.91 ;
        RECT 6.56 -0.085 6.89 0.855 ;
        RECT 4.295 -0.085 4.535 0.73 ;
        RECT 2.79 -0.085 3.12 0.485 ;
        RECT 0.805 -0.085 1.135 0.595 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.36 3.415 ;
        RECT 14.425 1.84 14.615 3.415 ;
        RECT 12.855 2.18 13.115 3.415 ;
        RECT 10.46 2.64 11.225 3.415 ;
        RECT 7.65 2.64 8.885 3.415 ;
        RECT 6.505 2.36 6.835 3.415 ;
        RECT 3.955 2.955 4.285 3.415 ;
        RECT 2.405 2.815 2.735 3.415 ;
        RECT 0.56 2.465 0.89 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 11.395 2.905 12.685 3.075 ;
      RECT 12.515 1.59 12.685 3.075 ;
      RECT 11.395 2.3 11.655 3.075 ;
      RECT 9.645 2.12 10.15 2.88 ;
      RECT 9.645 2.3 11.655 2.47 ;
      RECT 9.645 2.12 10.48 2.47 ;
      RECT 10.31 0.64 10.48 2.47 ;
      RECT 12.32 1.59 12.685 2.26 ;
      RECT 12.625 0.45 12.795 2.01 ;
      RECT 14.665 0.68 14.835 1.67 ;
      RECT 9.575 0.64 10.48 0.91 ;
      RECT 13.405 0.68 14.835 0.85 ;
      RECT 13.405 0.33 13.735 0.85 ;
      RECT 12.625 0.45 13.735 0.62 ;
      RECT 13.285 1.16 13.545 2.86 ;
      RECT 13.285 1.16 13.665 1.83 ;
      RECT 12.965 1.16 13.665 1.33 ;
      RECT 12.965 0.79 13.235 1.33 ;
      RECT 11.975 2.465 12.345 2.735 ;
      RECT 11.975 1.495 12.15 2.735 ;
      RECT 10.66 1.495 12.15 1.75 ;
      RECT 11.375 0.795 11.73 1.75 ;
      RECT 7.005 2.3 7.48 2.69 ;
      RECT 7.005 2.3 9.475 2.47 ;
      RECT 9.305 1.78 9.475 2.47 ;
      RECT 7.005 1.905 7.175 2.69 ;
      RECT 6.455 1.905 7.175 2.19 ;
      RECT 9.305 1.78 10.13 1.95 ;
      RECT 9.96 1.08 10.13 1.95 ;
      RECT 8.515 1.08 10.13 1.25 ;
      RECT 8.515 0.635 8.685 1.25 ;
      RECT 7.42 0.635 8.685 0.855 ;
      RECT 7.815 1.78 9.125 1.95 ;
      RECT 8.955 1.42 9.125 1.95 ;
      RECT 7.815 1.375 7.985 1.95 ;
      RECT 5.965 1.375 6.225 1.705 ;
      RECT 8.955 1.42 9.79 1.61 ;
      RECT 5.965 1.375 7.985 1.545 ;
      RECT 5.745 1.885 6.035 2.69 ;
      RECT 5.625 1.035 5.795 2.055 ;
      RECT 8.165 1.42 8.775 1.61 ;
      RECT 8.165 1.025 8.335 1.61 ;
      RECT 5.625 1.035 8.335 1.205 ;
      RECT 5.84 1.025 8.335 1.205 ;
      RECT 7.06 0.525 7.25 1.205 ;
      RECT 5.84 0.64 6.1 1.205 ;
      RECT 2.905 2.895 3.775 3.065 ;
      RECT 3.605 2.615 3.775 3.065 ;
      RECT 1.46 2.475 1.79 3.025 ;
      RECT 2.905 0.655 3.075 3.065 ;
      RECT 3.605 2.615 5.575 2.785 ;
      RECT 5.275 2.36 5.575 2.785 ;
      RECT 1.46 2.475 3.075 2.645 ;
      RECT 5.275 0.585 5.455 2.785 ;
      RECT 5.255 0.585 5.455 1.035 ;
      RECT 5.255 0.585 5.67 0.865 ;
      RECT 2.37 0.655 3.075 0.825 ;
      RECT 2.37 0.28 2.54 0.825 ;
      RECT 1.595 0.28 2.54 0.595 ;
      RECT 4.48 1.375 5.105 2.435 ;
      RECT 4.705 0.4 5.005 2.435 ;
      RECT 3.245 2.23 3.435 2.725 ;
      RECT 3.245 2.23 4.125 2.435 ;
      RECT 3.925 0.33 4.125 2.435 ;
      RECT 3.29 0.33 4.125 0.66 ;
      RECT 0.13 1.125 0.39 3.065 ;
      RECT 0.13 1.125 0.935 1.455 ;
      RECT 0.13 0.28 0.38 3.065 ;
      RECT 0.13 0.28 0.635 0.61 ;
  END
END scs130lp_sdfsbp_1

MACRO scs130lp_sdfsbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfsbp_2 0 0 ;
  SIZE 15.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.995 0.775 3.38 1.025 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.19 1.815 1.8 2.075 ;
        RECT 1.515 0.385 1.8 2.075 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8988 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.525 0.255 14.775 3.075 ;
        RECT 14.11 0.255 14.775 1.095 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.29 1.815 12.585 3.075 ;
        RECT 12.155 0.265 12.46 2.12 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.51 1.535 2.89 2.25 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.555 2.245 2.34 2.415 ;
        RECT 2.09 1.165 2.34 2.415 ;
        RECT 0.555 2.245 0.985 2.49 ;
        RECT 0.555 1.155 0.885 2.49 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
      ANTENNAGATEAREA 0.252 LAYER met1 ;
      ANTENNAMAXAREACAR 1.119048 LAYER li ;
      ANTENNAMAXAREACAR 1.119048 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.365079 LAYER li ;
      ANTENNAMAXSIDEAREACAR 1.365079 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.229365 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 10.655 1.92 10.945 2.15 ;
        RECT 7.295 1.965 10.945 2.105 ;
        RECT 7.295 1.92 7.585 2.15 ;
      LAYER li ;
        RECT 10.705 1.63 10.895 2.3 ;
        RECT 7.265 1.895 7.865 2.13 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.36 0.085 ;
        RECT 14.945 -0.085 15.215 1.095 ;
        RECT 13.655 -0.085 13.94 1.095 ;
        RECT 12.63 -0.085 12.965 1.105 ;
        RECT 11.55 -0.085 11.985 0.915 ;
        RECT 10.34 -0.085 10.67 0.915 ;
        RECT 8.14 -0.085 8.47 0.695 ;
        RECT 6.58 -0.085 6.91 0.97 ;
        RECT 4.145 -0.085 4.405 0.725 ;
        RECT 2.69 -0.085 3.02 0.535 ;
        RECT 0.83 -0.085 1.16 0.605 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.36 3.415 ;
        RECT 14.945 1.82 15.215 3.415 ;
        RECT 14.025 1.82 14.355 3.415 ;
        RECT 12.755 1.815 13.095 3.415 ;
        RECT 11.86 2.315 12.12 3.415 ;
        RECT 10.005 2.505 10.195 3.415 ;
        RECT 7.95 2.64 8.28 3.415 ;
        RECT 6.79 2.64 7.12 3.415 ;
        RECT 4.1 2.675 4.36 3.415 ;
        RECT 2.445 2.975 2.775 3.415 ;
        RECT 0.525 2.66 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 13.265 1.275 13.575 2.495 ;
      RECT 13.265 1.275 14.355 1.605 ;
      RECT 13.265 0.29 13.475 2.495 ;
      RECT 13.135 0.29 13.475 0.62 ;
      RECT 11.415 1.815 11.925 2.145 ;
      RECT 11.755 1.085 11.925 2.145 ;
      RECT 10.015 1.085 10.345 1.845 ;
      RECT 10.015 1.085 11.925 1.255 ;
      RECT 11.12 0.71 11.38 1.255 ;
      RECT 8.97 2.555 9.835 2.885 ;
      RECT 9.665 0.59 9.835 2.885 ;
      RECT 10.365 2.505 11.235 2.835 ;
      RECT 11.065 1.425 11.235 2.835 ;
      RECT 10.365 2.155 10.535 2.835 ;
      RECT 9.665 2.155 10.535 2.335 ;
      RECT 11.065 1.425 11.575 1.645 ;
      RECT 9.135 0.59 9.835 0.86 ;
      RECT 7.3 2.3 7.63 2.69 ;
      RECT 6.635 2.3 8.215 2.47 ;
      RECT 9.315 1.03 9.485 2.375 ;
      RECT 8.045 2.205 9.485 2.375 ;
      RECT 6.635 1.905 6.965 2.47 ;
      RECT 8.745 1.03 9.485 1.2 ;
      RECT 7.79 0.865 8.915 1.035 ;
      RECT 7.255 0.64 7.96 0.97 ;
      RECT 8.045 1.855 9.145 2.025 ;
      RECT 8.885 1.37 9.145 2.025 ;
      RECT 8.045 1.545 8.215 2.025 ;
      RECT 6.165 1.515 6.425 1.845 ;
      RECT 6.165 1.545 8.215 1.725 ;
      RECT 6.165 1.515 6.43 1.725 ;
      RECT 5.95 2.02 6.25 2.69 ;
      RECT 5.825 0.64 5.995 2.19 ;
      RECT 8.385 1.205 8.575 1.675 ;
      RECT 7.175 1.205 8.575 1.375 ;
      RECT 5.825 1.14 7.505 1.345 ;
      RECT 5.825 0.64 6.12 1.345 ;
      RECT 3.06 2.805 3.93 2.995 ;
      RECT 3.76 2.335 3.93 2.995 ;
      RECT 1.425 2.585 3.23 2.805 ;
      RECT 5.475 2.36 5.78 2.705 ;
      RECT 3.06 1.195 3.23 2.995 ;
      RECT 3.76 2.335 5.655 2.505 ;
      RECT 5.475 0.64 5.655 2.705 ;
      RECT 2.52 1.195 3.23 1.365 ;
      RECT 5.36 0.64 5.655 1.235 ;
      RECT 2.52 0.705 2.69 1.365 ;
      RECT 1.97 0.705 2.69 0.875 ;
      RECT 1.97 0.28 2.22 0.875 ;
      RECT 4.575 1.485 5.295 2.165 ;
      RECT 4.575 0.41 4.905 2.165 ;
      RECT 3.4 1.195 3.59 2.635 ;
      RECT 3.55 0.895 4.405 1.565 ;
      RECT 3.55 0.275 3.94 1.565 ;
      RECT 3.19 0.275 3.94 0.605 ;
      RECT 0.095 0.275 0.355 2.985 ;
      RECT 1.055 0.815 1.345 1.485 ;
      RECT 0.095 0.815 1.345 0.985 ;
      RECT 0.095 0.275 0.66 0.985 ;
  END
END scs130lp_sdfsbp_2

MACRO scs130lp_sdfsbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfsbp_lp 0 0 ;
  SIZE 16.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.215 1.45 4.645 1.78 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.46 2.3 1.79 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4026 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.615 1.85 16.21 2.89 ;
        RECT 16.04 0.35 16.21 2.89 ;
        RECT 15.88 0.35 16.21 0.81 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.995 1.61 14.245 3.02 ;
        RECT 13.565 0.265 14.075 0.725 ;
        RECT 13.565 1.61 14.245 1.78 ;
        RECT 13.565 0.265 13.795 1.78 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.365 1.11 3.685 1.78 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.51 1.11 2.835 1.79 ;
        RECT 1.565 1.11 2.835 1.28 ;
        RECT 0.93 0.855 2.275 1.185 ;
        RECT 1.565 0.81 2.275 1.28 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
      ANTENNAGATEAREA 0.626 LAYER met1 ;
      ANTENNAMAXAREACAR 0.401917 LAYER li ;
      ANTENNAMAXAREACAR 0.401917 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.453674 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.453674 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.092332 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 12.095 1.55 12.385 1.78 ;
        RECT 8.735 1.595 12.385 1.735 ;
        RECT 8.735 1.55 9.025 1.78 ;
      LAYER li ;
        RECT 11.985 1.55 12.355 1.89 ;
        RECT 8.795 1.55 9.065 1.88 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.32 0.245 ;
      LAYER li ;
        RECT 0 -0.085 16.32 0.085 ;
        RECT 15.09 -0.085 15.42 0.81 ;
        RECT 12.955 -0.085 13.285 0.725 ;
        RECT 11.59 -0.085 11.92 0.77 ;
        RECT 9.05 -0.085 9.38 1.02 ;
        RECT 7.315 -0.085 7.565 0.695 ;
        RECT 4.655 -0.085 4.825 0.92 ;
        RECT 2.995 -0.085 3.325 0.58 ;
        RECT 1.055 -0.085 1.385 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.32 3.575 ;
      LAYER li ;
        RECT 0 3.245 16.32 3.415 ;
        RECT 15.085 1.85 15.415 3.415 ;
        RECT 13.545 1.98 13.795 3.415 ;
        RECT 11.51 2.465 11.84 3.415 ;
        RECT 8.8 2.865 9.13 3.415 ;
        RECT 7.74 2.865 8.07 3.415 ;
        RECT 4.38 2.31 4.71 3.415 ;
        RECT 2.755 2.67 3.085 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 14.46 1.49 14.885 2.89 ;
      RECT 14.46 1.49 15.725 1.66 ;
      RECT 15.395 0.99 15.725 1.66 ;
      RECT 14.46 0.35 14.63 2.89 ;
      RECT 14.3 0.35 14.63 0.81 ;
      RECT 12.21 2.895 13.365 3.065 ;
      RECT 13.195 1.17 13.365 3.065 ;
      RECT 10.205 2.075 10.535 3.065 ;
      RECT 12.21 2.075 12.46 3.065 ;
      RECT 10.205 2.115 12.46 2.285 ;
      RECT 11.16 0.95 11.33 2.285 ;
      RECT 12.99 1.17 13.365 1.84 ;
      RECT 10.325 0.95 11.33 1.12 ;
      RECT 10.325 0.31 10.655 1.12 ;
      RECT 12.64 2.02 13.015 2.715 ;
      RECT 12.64 1.2 12.81 2.715 ;
      RECT 11.51 1.2 11.775 1.885 ;
      RECT 11.51 1.2 12.81 1.37 ;
      RECT 12.165 0.265 12.495 1.37 ;
      RECT 4.91 2.895 7.56 3.065 ;
      RECT 7.39 2.515 7.56 3.065 ;
      RECT 5.96 1.3 6.13 3.065 ;
      RECT 4.91 2.31 5.24 3.065 ;
      RECT 7.39 2.515 9.985 2.685 ;
      RECT 9.815 1.155 9.985 2.685 ;
      RECT 10.715 1.605 10.98 1.935 ;
      RECT 5.67 1.3 6.13 1.78 ;
      RECT 9.815 1.605 10.98 1.775 ;
      RECT 5.67 1.3 6.905 1.63 ;
      RECT 9.815 1.155 10.145 1.775 ;
      RECT 5.67 0.615 5.84 1.78 ;
      RECT 5.365 0.615 5.84 1.005 ;
      RECT 6.31 2.075 6.64 2.715 ;
      RECT 6.31 2.075 7.255 2.245 ;
      RECT 7.085 0.875 7.255 2.245 ;
      RECT 8.005 1.575 8.615 1.905 ;
      RECT 8.445 1.2 8.615 1.905 ;
      RECT 9.275 1.2 9.605 1.87 ;
      RECT 8.445 1.2 9.605 1.37 ;
      RECT 8.7 0.265 8.87 1.37 ;
      RECT 6.45 0.605 6.78 1.065 ;
      RECT 6.45 0.875 7.915 1.045 ;
      RECT 7.745 0.265 7.915 1.045 ;
      RECT 7.745 0.265 8.87 0.435 ;
      RECT 7.435 2.085 8.6 2.335 ;
      RECT 7.435 1.225 7.765 2.335 ;
      RECT 7.435 1.225 8.265 1.395 ;
      RECT 8.095 0.615 8.265 1.395 ;
      RECT 8.095 0.615 8.52 1.02 ;
      RECT 5.45 1.96 5.78 2.715 ;
      RECT 1.735 1.97 2.065 2.715 ;
      RECT 1.735 1.97 3.185 2.14 ;
      RECT 3.015 0.76 3.185 2.14 ;
      RECT 5.32 1.185 5.49 2.13 ;
      RECT 5.015 1.185 5.49 1.355 ;
      RECT 4.295 1.1 5.185 1.27 ;
      RECT 5.015 0.265 5.185 1.355 ;
      RECT 4.295 0.265 4.465 1.27 ;
      RECT 2.455 0.76 3.675 0.93 ;
      RECT 3.505 0.265 3.675 0.93 ;
      RECT 6.02 0.265 6.27 0.855 ;
      RECT 2.455 0.265 2.625 0.93 ;
      RECT 2.175 0.265 2.625 0.63 ;
      RECT 5.015 0.265 6.27 0.435 ;
      RECT 3.505 0.265 4.465 0.435 ;
      RECT 3.85 1.96 4.18 3.065 ;
      RECT 3.85 1.96 5.14 2.13 ;
      RECT 4.825 1.555 5.14 2.13 ;
      RECT 3.865 0.615 4.035 3.065 ;
      RECT 3.865 0.615 4.115 1.005 ;
      RECT 3.285 2.32 3.615 3.065 ;
      RECT 1.205 2.895 2.575 3.065 ;
      RECT 2.405 2.32 2.575 3.065 ;
      RECT 1.205 2.025 1.535 3.065 ;
      RECT 2.405 2.32 3.615 2.49 ;
      RECT 0.115 0.265 0.445 3.065 ;
      RECT 0.115 1.425 1.385 1.755 ;
      RECT 0.115 0.265 0.565 1.755 ;
  END
END scs130lp_sdfsbp_lp

MACRO scs130lp_sdfstp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfstp_1 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.95 0.78 4.285 1.825 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.015 1.53 2.255 1.84 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.035 1.85 14.315 3.075 ;
        RECT 14.065 0.325 14.315 3.075 ;
        RECT 13.925 0.325 14.315 1.125 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.155 1.17 0.62 1.84 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.43 0.265 3.275 0.64 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.45 1.585 11.66 1.765 ;
        RECT 10.45 0.265 10.62 1.765 ;
        RECT 7.835 0.265 10.62 0.64 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 14.4 0.085 ;
        RECT 13.4 -0.085 13.755 1.125 ;
        RECT 11.495 -0.085 11.825 0.995 ;
        RECT 7.485 0.82 8.855 1.01 ;
        RECT 7.485 -0.085 7.655 1.01 ;
        RECT 6.44 -0.085 6.77 0.665 ;
        RECT 3.95 -0.085 4.2 0.61 ;
        RECT 1.745 -0.085 2.015 1.015 ;
        RECT 0.165 -0.085 0.495 1 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 14.4 3.415 ;
        RECT 13.425 1.815 13.865 3.415 ;
        RECT 12.01 2.465 12.34 3.415 ;
        RECT 11.09 2.465 11.35 3.415 ;
        RECT 7.97 2.155 8.31 3.415 ;
        RECT 6.44 2.37 6.72 3.415 ;
        RECT 4.24 2.845 4.57 3.415 ;
        RECT 2.375 2.81 2.705 3.415 ;
        RECT 0.56 2.35 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 12.95 1.295 13.255 2.495 ;
      RECT 12.95 1.295 13.895 1.625 ;
      RECT 12.95 0.81 13.23 2.495 ;
      RECT 12.51 1.235 12.77 2.795 ;
      RECT 10.79 1.235 12.77 1.415 ;
      RECT 11.995 0.665 12.325 1.415 ;
      RECT 11.52 1.935 11.76 2.795 ;
      RECT 11.52 1.935 12.34 2.255 ;
      RECT 12.09 1.585 12.34 2.255 ;
      RECT 9.64 1.935 12.34 2.115 ;
      RECT 9.64 0.81 10.28 2.115 ;
      RECT 9.01 2.795 10.92 2.965 ;
      RECT 10.63 2.465 10.92 2.965 ;
      RECT 9.01 2.625 9.34 2.965 ;
      RECT 8.49 2.155 8.82 2.755 ;
      RECT 10.08 2.285 10.41 2.625 ;
      RECT 8.49 2.285 10.41 2.455 ;
      RECT 4.74 2.865 6.25 3.035 ;
      RECT 6.08 1.595 6.25 3.035 ;
      RECT 6.89 2.84 7.8 3.01 ;
      RECT 7.63 1.815 7.8 3.01 ;
      RECT 4.74 2.695 5 3.035 ;
      RECT 6.89 1.945 7.06 3.01 ;
      RECT 6.08 1.945 7.06 2.115 ;
      RECT 9.14 1.815 9.47 2.105 ;
      RECT 7.63 1.815 9.47 1.985 ;
      RECT 6.08 1.595 6.41 2.115 ;
      RECT 5.72 0.325 5.9 2.69 ;
      RECT 8.365 1.245 8.695 1.645 ;
      RECT 5.72 1.245 8.695 1.425 ;
      RECT 5.72 0.325 5.92 0.725 ;
      RECT 7.23 1.595 7.46 2.67 ;
      RECT 6.62 1.595 7.46 1.775 ;
      RECT 6.47 0.835 7.315 1.075 ;
      RECT 7.055 0.66 7.315 1.075 ;
      RECT 5.37 0.265 5.55 1.845 ;
      RECT 4.37 0.265 4.66 0.61 ;
      RECT 4.37 0.265 5.55 0.435 ;
      RECT 2.885 2.895 4.06 3.065 ;
      RECT 3.89 2.495 4.06 3.065 ;
      RECT 2.885 2.45 3.055 3.065 ;
      RECT 5.2 2.295 5.55 2.69 ;
      RECT 3.89 2.495 4.57 2.665 ;
      RECT 1.37 2.45 3.055 2.64 ;
      RECT 5.03 0.605 5.2 2.525 ;
      RECT 4.4 2.355 5.55 2.525 ;
      RECT 2.425 1.19 2.595 2.64 ;
      RECT 1.37 2.35 1.7 2.64 ;
      RECT 0.955 1.19 2.595 1.36 ;
      RECT 0.955 0.685 1.285 1.36 ;
      RECT 4.87 0.605 5.2 0.805 ;
      RECT 3.61 1.995 4.025 2.315 ;
      RECT 3.61 1.995 4.835 2.185 ;
      RECT 3.61 0.28 3.78 2.315 ;
      RECT 3.47 0.28 3.78 0.61 ;
      RECT 3.225 1.62 3.44 2.725 ;
      RECT 2.765 1.62 3.44 1.79 ;
      RECT 2.765 0.81 3.025 1.79 ;
      RECT 2.215 0.81 3.025 1.02 ;
      RECT 0.095 2.01 0.39 2.7 ;
      RECT 1.855 2.01 2.185 2.28 ;
      RECT 0.095 2.01 2.185 2.18 ;
  END
END scs130lp_sdfstp_1

MACRO scs130lp_sdfstp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfstp_2 0 0 ;
  SIZE 15.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.305 0.78 4.685 1.825 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.95 2.255 2.225 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.555 0.965 15.275 1.995 ;
        RECT 14.39 1.825 14.59 3.075 ;
        RECT 14.39 0.255 14.59 1.135 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.15 0.55 1.78 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 0.265 3.765 1.38 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.87 1.585 12.09 1.765 ;
        RECT 10.87 0.265 11.04 1.765 ;
        RECT 8.315 0.265 11.04 0.5 ;
        RECT 8.315 0.265 9.925 0.64 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.36 0.085 ;
        RECT 14.76 -0.085 15.09 0.795 ;
        RECT 13.84 -0.085 14.17 1.095 ;
        RECT 11.885 -0.085 12.215 0.995 ;
        RECT 7.965 0.81 9.54 1.01 ;
        RECT 7.965 -0.085 8.135 1.01 ;
        RECT 6.95 -0.085 7.28 0.555 ;
        RECT 4.4 -0.085 4.655 0.61 ;
        RECT 1.985 -0.085 2.62 0.98 ;
        RECT 0.405 -0.085 0.735 0.98 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.36 3.415 ;
        RECT 14.76 2.165 15.09 3.415 ;
        RECT 13.855 1.825 14.22 3.415 ;
        RECT 12.44 2.46 12.76 3.415 ;
        RECT 11.53 2.275 11.785 3.415 ;
        RECT 8.52 2.075 8.745 3.415 ;
        RECT 6.98 2.275 7.31 3.415 ;
        RECT 4.5 2.835 4.83 3.415 ;
        RECT 2.765 2.3 3.025 3.415 ;
        RECT 0.585 2.815 0.915 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 13.39 1.315 13.685 2.485 ;
      RECT 13.39 1.315 14.335 1.645 ;
      RECT 13.39 0.7 13.67 2.485 ;
      RECT 12.93 1.235 13.2 2.79 ;
      RECT 11.22 1.235 13.2 1.415 ;
      RECT 12.425 0.665 12.755 1.415 ;
      RECT 11.955 1.935 12.25 2.55 ;
      RECT 11.955 1.935 12.76 2.255 ;
      RECT 12.5 1.585 12.76 2.255 ;
      RECT 10.08 1.935 12.76 2.105 ;
      RECT 10.08 1.915 10.7 2.105 ;
      RECT 10.095 0.67 10.7 2.105 ;
      RECT 9.42 2.795 11.36 2.965 ;
      RECT 11.06 2.275 11.36 2.965 ;
      RECT 9.42 2.615 9.75 2.965 ;
      RECT 8.915 2.075 9.21 2.755 ;
      RECT 10.51 2.275 10.84 2.615 ;
      RECT 8.915 2.275 10.84 2.445 ;
      RECT 5 2.705 6.79 3.035 ;
      RECT 6.62 1.935 6.79 3.035 ;
      RECT 7.48 2.565 8.35 2.735 ;
      RECT 8.18 1.735 8.35 2.735 ;
      RECT 5.91 1.375 6.09 3.035 ;
      RECT 7.48 1.935 7.65 2.735 ;
      RECT 6.62 1.935 7.65 2.105 ;
      RECT 9.61 1.735 9.91 2.095 ;
      RECT 8.18 1.735 9.91 1.905 ;
      RECT 5.88 0.255 6.07 1.705 ;
      RECT 4.825 0.255 5.12 0.61 ;
      RECT 4.825 0.255 6.07 0.425 ;
      RECT 6.26 1.225 6.45 2.385 ;
      RECT 6.26 1.225 9.085 1.415 ;
      RECT 6.26 0.325 6.43 2.385 ;
      RECT 6.24 0.325 6.43 0.715 ;
      RECT 7.82 1.585 8.01 2.385 ;
      RECT 6.845 1.585 8.01 1.765 ;
      RECT 1.43 2.815 2.595 3.075 ;
      RECT 2.425 1.15 2.595 3.075 ;
      RECT 3.195 2.8 4.32 2.97 ;
      RECT 4.15 2.495 4.32 2.97 ;
      RECT 3.195 1.95 3.365 2.97 ;
      RECT 4.15 2.495 4.83 2.665 ;
      RECT 5.38 2.185 5.74 2.525 ;
      RECT 4.66 2.355 5.74 2.525 ;
      RECT 5.38 0.595 5.71 2.525 ;
      RECT 2.425 1.95 3.365 2.12 ;
      RECT 1.195 1.15 2.595 1.405 ;
      RECT 1.195 0.65 1.525 1.405 ;
      RECT 3.965 1.995 4.305 2.325 ;
      RECT 3.965 1.995 5.135 2.185 ;
      RECT 4.855 1.245 5.135 2.185 ;
      RECT 3.965 0.28 4.135 2.325 ;
      RECT 3.965 0.28 4.23 0.61 ;
      RECT 3.535 1.55 3.785 2.63 ;
      RECT 2.79 1.55 3.785 1.78 ;
      RECT 2.79 0.65 3.085 1.78 ;
      RECT 0.155 2.395 0.415 3.065 ;
      RECT 0.155 2.395 2.245 2.645 ;
      RECT 6.825 0.725 7.795 1.055 ;
  END
END scs130lp_sdfstp_2

MACRO scs130lp_sdfstp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfstp_4 0 0 ;
  SIZE 15.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.205 0.83 4.78 1.775 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.935 2.255 2.155 ;
        RECT 0.72 1.87 2.255 2.155 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.07 1.765 15.685 1.935 ;
        RECT 15.035 1.075 15.685 1.935 ;
        RECT 14.97 1.765 15.16 3.075 ;
        RECT 14.94 0.255 15.13 1.255 ;
        RECT 14.08 1.075 15.685 1.255 ;
        RECT 14.07 1.765 14.3 3.075 ;
        RECT 14.08 0.255 14.27 1.255 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.14 0.55 1.765 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.435 0.39 3.695 1.76 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.685 1.585 11.895 1.765 ;
        RECT 10.685 0.255 10.855 1.765 ;
        RECT 8.305 0.255 10.855 0.665 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.84 0.085 ;
        RECT 15.3 -0.085 15.63 0.905 ;
        RECT 14.44 -0.085 14.77 0.905 ;
        RECT 13.58 -0.085 13.91 1.13 ;
        RECT 11.745 -0.085 12.075 1.005 ;
        RECT 7.965 0.835 9.315 1.185 ;
        RECT 7.965 -0.085 8.135 1.185 ;
        RECT 6.91 -0.085 7.24 0.78 ;
        RECT 4.41 -0.085 4.66 0.66 ;
        RECT 1.855 -0.085 2.185 0.97 ;
        RECT 0.275 -0.085 0.605 0.97 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.84 3.415 ;
        RECT 15.33 2.105 15.66 3.415 ;
        RECT 14.47 2.105 14.8 3.415 ;
        RECT 13.65 1.815 13.9 3.415 ;
        RECT 12.23 2.46 12.525 3.415 ;
        RECT 11.34 2.63 11.55 3.415 ;
        RECT 8.3 2.135 8.63 3.415 ;
        RECT 6.89 2.435 7.08 3.415 ;
        RECT 4.35 2.795 4.61 3.415 ;
        RECT 2.645 2.725 2.855 3.415 ;
        RECT 0.525 2.665 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 13.16 1.425 13.48 3.075 ;
      RECT 13.16 1.425 14.855 1.595 ;
      RECT 13.16 0.255 13.41 3.075 ;
      RECT 12.695 1.235 12.99 2.79 ;
      RECT 11.025 1.235 12.99 1.415 ;
      RECT 11.025 1.175 12.56 1.415 ;
      RECT 12.265 0.675 12.56 1.415 ;
      RECT 11.77 1.935 12.06 2.96 ;
      RECT 11.77 1.935 12.465 2.255 ;
      RECT 12.11 1.585 12.465 2.255 ;
      RECT 9.87 1.935 12.465 2.125 ;
      RECT 9.87 0.835 10.515 2.125 ;
      RECT 9.25 2.695 11.12 3.025 ;
      RECT 9.25 2.645 9.58 3.025 ;
      RECT 8.8 2.295 9 2.635 ;
      RECT 10.3 2.295 10.63 2.525 ;
      RECT 8.8 2.295 10.63 2.475 ;
      RECT 4.78 2.805 6.72 3.075 ;
      RECT 6.54 2.095 6.72 3.075 ;
      RECT 7.25 2.785 8.12 2.955 ;
      RECT 7.95 1.795 8.12 2.955 ;
      RECT 4.78 2.795 5.93 3.075 ;
      RECT 5.76 1.295 5.93 3.075 ;
      RECT 7.25 2.095 7.42 2.955 ;
      RECT 6.54 2.095 7.42 2.265 ;
      RECT 9.36 1.795 9.69 2.015 ;
      RECT 7.95 1.795 9.69 1.965 ;
      RECT 5.85 0.255 6.02 1.965 ;
      RECT 4.83 0.255 5.07 0.66 ;
      RECT 4.83 0.255 6.02 0.425 ;
      RECT 6.1 2.305 6.37 2.635 ;
      RECT 6.19 0.535 6.37 2.635 ;
      RECT 8.605 1.355 8.935 1.625 ;
      RECT 6.19 1.355 8.935 1.545 ;
      RECT 6.19 0.535 6.45 0.865 ;
      RECT 6.785 0.95 7.785 1.185 ;
      RECT 7.595 0.735 7.785 1.185 ;
      RECT 7.59 1.715 7.78 2.615 ;
      RECT 6.695 1.715 7.78 1.925 ;
      RECT 3.025 2.905 4.18 3.075 ;
      RECT 3.955 2.455 4.18 3.075 ;
      RECT 1.37 2.905 2.475 3.075 ;
      RECT 3.025 2.385 3.195 3.075 ;
      RECT 2.305 2.385 2.475 3.075 ;
      RECT 1.37 2.665 1.7 3.075 ;
      RECT 3.955 2.455 5.59 2.625 ;
      RECT 5.34 0.595 5.59 2.625 ;
      RECT 2.305 2.385 3.195 2.555 ;
      RECT 2.425 1.215 2.595 2.555 ;
      RECT 1.065 1.215 2.595 1.54 ;
      RECT 1.065 0.64 1.395 1.54 ;
      RECT 5.34 0.595 5.68 0.805 ;
      RECT 3.825 2.025 4.985 2.285 ;
      RECT 3.865 1.945 4.985 2.285 ;
      RECT 3.865 0.33 4.035 2.285 ;
      RECT 3.865 0.33 4.24 0.66 ;
      RECT 3.365 1.93 3.625 2.735 ;
      RECT 2.765 1.93 3.625 2.1 ;
      RECT 2.765 0.64 3.025 2.1 ;
      RECT 2.355 0.64 3.025 0.97 ;
      RECT 0.095 2.325 0.355 3.045 ;
      RECT 1.87 2.325 2.135 2.735 ;
      RECT 0.095 2.325 2.135 2.495 ;
  END
END scs130lp_sdfstp_4

MACRO scs130lp_sdfstp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfstp_lp 0 0 ;
  SIZE 15.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.215 1.51 4.645 1.84 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.46 2.3 1.79 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.205 1.85 15.725 2.89 ;
        RECT 15.485 0.265 15.725 2.89 ;
        RECT 15.395 0.265 15.725 0.725 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.365 1.16 3.685 1.83 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.51 1.11 2.835 1.79 ;
        RECT 1.565 1.11 2.835 1.28 ;
        RECT 0.75 0.855 2.275 1.185 ;
        RECT 1.565 0.81 2.275 1.28 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
      ANTENNAGATEAREA 0.626 LAYER met1 ;
      ANTENNAMAXAREACAR 0.933067 LAYER li ;
      ANTENNAMAXAREACAR 0.933067 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.776358 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.776358 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.092332 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 12.095 1.92 12.385 2.15 ;
        RECT 8.735 1.965 12.385 2.105 ;
        RECT 8.735 1.92 9.025 2.15 ;
      LAYER li ;
        RECT 12.1 1.265 12.43 2.15 ;
        RECT 8.795 1.605 9.1 2.15 ;
    END
  END SETB
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.84 0.085 ;
        RECT 14.605 -0.085 14.935 0.725 ;
        RECT 13.255 -0.085 13.585 0.725 ;
        RECT 11.375 -0.085 11.705 0.735 ;
        RECT 9.085 -0.085 9.415 1.065 ;
        RECT 7.315 -0.085 7.565 0.685 ;
        RECT 4.63 -0.085 4.8 0.98 ;
        RECT 3.025 -0.085 3.275 0.58 ;
        RECT 1.055 -0.085 1.385 0.675 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.84 3.415 ;
        RECT 14.675 1.85 15.005 3.415 ;
        RECT 13.665 1.755 13.915 3.415 ;
        RECT 11.545 2.68 11.875 3.415 ;
        RECT 8.79 2.855 9.12 3.415 ;
        RECT 7.44 2.855 7.77 3.415 ;
        RECT 4.375 2.37 4.705 3.415 ;
        RECT 2.755 2.67 3.085 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 14.095 0.99 14.475 2.89 ;
      RECT 14.91 0.99 15.24 1.66 ;
      RECT 14.095 0.99 15.24 1.16 ;
      RECT 14.095 0.265 14.265 2.89 ;
      RECT 13.815 0.265 14.265 0.725 ;
      RECT 12.325 2.895 13.485 3.065 ;
      RECT 13.315 0.905 13.485 3.065 ;
      RECT 10.24 2.075 10.57 3.065 ;
      RECT 12.325 2.33 12.655 3.065 ;
      RECT 10.24 2.33 12.655 2.5 ;
      RECT 11.235 0.915 11.405 2.5 ;
      RECT 13.315 0.905 13.645 1.575 ;
      RECT 10.085 0.915 11.405 1.085 ;
      RECT 10.085 0.31 10.53 1.085 ;
      RECT 12.885 0.915 13.135 2.715 ;
      RECT 11.585 0.915 11.89 1.885 ;
      RECT 11.585 0.915 13.135 1.085 ;
      RECT 12.465 0.265 12.795 1.085 ;
      RECT 4.905 2.895 6.98 3.065 ;
      RECT 6.81 2.505 6.98 3.065 ;
      RECT 5.95 1.3 6.12 3.065 ;
      RECT 4.905 2.37 5.235 3.065 ;
      RECT 6.81 2.505 10.02 2.675 ;
      RECT 9.85 1.3 10.02 2.675 ;
      RECT 10.75 1.46 11.055 1.935 ;
      RECT 5.63 1.3 6.12 1.84 ;
      RECT 9.85 1.46 11.055 1.63 ;
      RECT 5.63 1.3 6.895 1.63 ;
      RECT 9.85 1.3 10.18 1.63 ;
      RECT 5.63 0.615 5.8 1.84 ;
      RECT 5.34 0.615 5.8 0.98 ;
      RECT 6.3 2.075 6.63 2.715 ;
      RECT 6.3 2.075 7.245 2.245 ;
      RECT 7.075 0.865 7.245 2.245 ;
      RECT 9.31 1.245 9.64 1.915 ;
      RECT 7.995 1.565 8.615 1.895 ;
      RECT 8.445 1.245 8.615 1.895 ;
      RECT 8.445 1.245 9.64 1.415 ;
      RECT 8.735 0.265 8.905 1.415 ;
      RECT 6.395 0.865 7.245 1.065 ;
      RECT 6.395 0.865 7.915 1.035 ;
      RECT 7.745 0.265 7.915 1.035 ;
      RECT 6.395 0.605 6.725 1.065 ;
      RECT 7.745 0.265 8.905 0.435 ;
      RECT 7.425 2.075 8.59 2.325 ;
      RECT 7.425 1.215 7.755 2.325 ;
      RECT 7.425 1.215 8.265 1.385 ;
      RECT 8.095 0.615 8.265 1.385 ;
      RECT 8.095 0.615 8.555 1.065 ;
      RECT 5.44 2.02 5.77 2.715 ;
      RECT 1.735 1.97 2.065 2.715 ;
      RECT 5.28 1.16 5.45 2.19 ;
      RECT 1.735 1.97 3.185 2.14 ;
      RECT 3.015 0.76 3.185 2.14 ;
      RECT 4.24 1.16 5.45 1.33 ;
      RECT 4.99 0.265 5.16 1.33 ;
      RECT 4.24 0.265 4.41 1.33 ;
      RECT 5.98 0.265 6.15 1.065 ;
      RECT 2.455 0.76 3.625 0.93 ;
      RECT 3.455 0.265 3.625 0.93 ;
      RECT 2.455 0.265 2.625 0.93 ;
      RECT 2.205 0.265 2.625 0.63 ;
      RECT 4.99 0.265 6.15 0.435 ;
      RECT 3.455 0.265 4.41 0.435 ;
      RECT 3.845 2.02 4.175 3.065 ;
      RECT 3.845 2.02 5.1 2.19 ;
      RECT 4.825 1.555 5.1 2.19 ;
      RECT 3.865 0.615 4.035 3.065 ;
      RECT 3.81 0.615 4.06 0.98 ;
      RECT 1.205 2.895 2.415 3.065 ;
      RECT 2.245 2.32 2.415 3.065 ;
      RECT 3.365 2.01 3.615 3.05 ;
      RECT 1.205 2.01 1.535 3.065 ;
      RECT 2.245 2.32 3.615 2.49 ;
      RECT 0.115 0.265 0.445 3.065 ;
      RECT 0.115 1.46 1.385 1.79 ;
      RECT 0.115 0.265 0.595 0.675 ;
  END
END scs130lp_sdfstp_lp

MACRO scs130lp_sdfxbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfxbp_1 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.825 1.12 8.52 1.455 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.02 1.345 1.52 2.12 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.99 1.345 13.405 2.145 ;
        RECT 12.99 0.375 13.285 2.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6153 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.045 0.375 14.315 3.075 ;
        RECT 13.845 0.375 14.315 1.175 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.14 0.55 2.12 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.975 0.265 3.215 1.39 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 14.4 0.085 ;
        RECT 13.455 -0.085 13.675 1.175 ;
        RECT 11.98 -0.085 12.27 0.805 ;
        RECT 10.68 -0.085 11.01 1.215 ;
        RECT 7.805 -0.085 8.08 0.95 ;
        RECT 4.575 -0.085 4.905 1.165 ;
        RECT 1.855 -0.085 2.185 0.835 ;
        RECT 0.165 -0.085 0.495 0.97 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 14.4 3.415 ;
        RECT 13.545 2.665 13.875 3.415 ;
        RECT 12.53 2.665 12.86 3.415 ;
        RECT 10.98 2.145 11.335 3.415 ;
        RECT 7.83 2.685 8.16 3.415 ;
        RECT 4.32 2.725 4.65 3.415 ;
        RECT 3.315 2.725 3.575 3.415 ;
        RECT 0.525 2.63 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 12.005 2.325 13.875 2.495 ;
      RECT 13.625 1.345 13.875 2.495 ;
      RECT 12.005 1.815 12.81 2.495 ;
      RECT 12.64 0.475 12.81 2.495 ;
      RECT 12.44 0.475 12.81 0.805 ;
      RECT 11.505 0.975 11.785 2.755 ;
      RECT 10.41 1.805 11.785 1.975 ;
      RECT 10.41 1.785 10.74 1.975 ;
      RECT 11.505 0.975 12.46 1.645 ;
      RECT 11.18 0.595 11.685 1.265 ;
      RECT 9.53 1.445 9.86 2.175 ;
      RECT 11.005 1.445 11.335 1.635 ;
      RECT 9.53 1.445 11.335 1.615 ;
      RECT 9.745 0.795 10.075 1.615 ;
      RECT 8.91 2.725 10.81 2.945 ;
      RECT 10.48 2.245 10.81 2.945 ;
      RECT 8.91 2.685 9.24 2.945 ;
      RECT 10.02 2.345 10.24 2.555 ;
      RECT 10.03 1.875 10.24 2.555 ;
      RECT 6.565 2.345 10.24 2.515 ;
      RECT 9.085 0.67 9.255 2.515 ;
      RECT 6.565 1.685 6.735 2.515 ;
      RECT 3.795 1.685 5.05 2.215 ;
      RECT 3.795 1.685 6.735 1.855 ;
      RECT 3.795 0.615 4.065 2.215 ;
      RECT 9.085 0.67 9.575 1 ;
      RECT 8.32 1.625 8.915 2.175 ;
      RECT 8.69 0.615 8.915 2.175 ;
      RECT 7.405 1.625 8.915 1.795 ;
      RECT 7.405 1.125 7.655 1.795 ;
      RECT 8.25 0.615 8.915 0.945 ;
      RECT 6.905 1.975 7.635 2.165 ;
      RECT 6.905 0.615 7.165 2.165 ;
      RECT 6.905 0.615 7.635 0.945 ;
      RECT 6.95 0.255 7.28 0.945 ;
      RECT 4.94 2.895 6.895 3.065 ;
      RECT 6.565 2.685 6.895 3.065 ;
      RECT 4.94 2.725 5.27 3.065 ;
      RECT 5.5 0.255 5.795 0.98 ;
      RECT 6.38 0.255 6.71 0.855 ;
      RECT 5.5 0.255 6.71 0.435 ;
      RECT 6.055 2.025 6.385 2.725 ;
      RECT 5.39 2.025 6.385 2.215 ;
      RECT 1.315 2.895 3.145 3.065 ;
      RECT 2.975 1.56 3.145 3.065 ;
      RECT 1.315 2.835 2.425 3.065 ;
      RECT 2.255 1.205 2.425 3.065 ;
      RECT 5.545 2.385 5.875 2.725 ;
      RECT 2.975 2.385 5.875 2.555 ;
      RECT 2.975 1.56 3.555 1.73 ;
      RECT 3.385 0.265 3.555 1.73 ;
      RECT 4.235 1.335 6.2 1.505 ;
      RECT 5.965 0.65 6.2 1.505 ;
      RECT 1.7 1.205 2.425 1.415 ;
      RECT 4.235 0.265 4.405 1.505 ;
      RECT 1.7 1.005 1.87 1.415 ;
      RECT 1.01 1.005 1.87 1.175 ;
      RECT 1.01 0.64 1.34 1.175 ;
      RECT 3.385 0.265 4.405 0.435 ;
      RECT 2.595 0.64 2.805 2.725 ;
      RECT 2.355 0.64 2.805 0.97 ;
      RECT 0.095 2.29 0.355 3.065 ;
      RECT 1.745 2.29 2.075 2.665 ;
      RECT 0.095 2.29 2.075 2.46 ;
  END
END scs130lp_sdfxbp_1

MACRO scs130lp_sdfxbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfxbp_2 0 0 ;
  SIZE 15.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.345 1.14 8.55 1.395 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.04 1.385 1.85 2.12 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.11 1.875 12.92 2.205 ;
        RECT 12.11 1.05 12.87 1.22 ;
        RECT 12.64 0.26 12.87 1.22 ;
        RECT 12.11 1.05 12.335 2.205 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.555 0.255 14.815 3.075 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.185 0.805 2.12 ;
        RECT 0.085 1.145 0.755 2.12 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.02 0.265 3.285 1.485 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.36 0.085 ;
        RECT 14.985 -0.085 15.255 1.09 ;
        RECT 14.045 -0.085 14.375 0.885 ;
        RECT 13.04 -0.085 13.385 1.14 ;
        RECT 12.14 -0.085 12.47 0.88 ;
        RECT 11.01 -0.085 11.34 1.21 ;
        RECT 7.93 -0.085 8.18 0.97 ;
        RECT 4.71 -0.085 5.04 1.165 ;
        RECT 1.785 -0.085 2.115 0.86 ;
        RECT 0.095 -0.085 0.425 0.975 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.36 3.415 ;
        RECT 14.985 1.815 15.255 3.415 ;
        RECT 14.125 2.105 14.335 3.415 ;
        RECT 13.02 2.715 13.35 3.415 ;
        RECT 12.16 2.715 12.49 3.415 ;
        RECT 10.915 2.145 11.39 3.415 ;
        RECT 7.81 2.705 8.14 3.415 ;
        RECT 4.415 2.715 4.745 3.415 ;
        RECT 3.36 2.715 3.61 3.415 ;
        RECT 0.595 2.63 0.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 13.545 1.755 13.875 2.485 ;
      RECT 13.545 1.755 14.375 1.925 ;
      RECT 14.025 1.055 14.375 1.925 ;
      RECT 13.555 1.055 14.375 1.225 ;
      RECT 13.555 0.325 13.855 1.225 ;
      RECT 11.56 1.795 11.94 2.755 ;
      RECT 11.69 0.59 11.94 2.755 ;
      RECT 11.56 2.375 13.32 2.545 ;
      RECT 13.15 1.405 13.32 2.545 ;
      RECT 10.61 1.795 11.94 1.975 ;
      RECT 10.61 1.72 10.94 1.975 ;
      RECT 12.505 1.405 13.32 1.655 ;
      RECT 12.505 1.405 13.855 1.585 ;
      RECT 11.52 0.59 11.94 1.21 ;
      RECT 10.045 0.66 10.36 2.775 ;
      RECT 11.18 1.38 11.51 1.625 ;
      RECT 10.045 1.38 11.51 1.55 ;
      RECT 9.615 0.66 9.875 2.775 ;
      RECT 6.625 2.365 9.875 2.535 ;
      RECT 6.625 1.675 6.795 2.535 ;
      RECT 3.87 2.035 5.145 2.205 ;
      RECT 4.815 1.675 5.145 2.205 ;
      RECT 3.87 0.635 4.2 2.205 ;
      RECT 4.815 1.675 6.795 1.845 ;
      RECT 8.32 1.565 8.65 2.195 ;
      RECT 7.59 1.565 8.65 1.77 ;
      RECT 7.59 1.565 9.05 1.735 ;
      RECT 8.72 0.64 9.05 1.735 ;
      RECT 8.35 0.64 9.05 0.97 ;
      RECT 6.995 1.94 7.515 2.195 ;
      RECT 6.995 0.255 7.175 2.195 ;
      RECT 6.995 0.64 7.76 0.97 ;
      RECT 6.995 0.255 7.395 0.97 ;
      RECT 5.035 2.905 6.955 3.075 ;
      RECT 6.625 2.705 6.955 3.075 ;
      RECT 5.035 2.715 5.365 3.075 ;
      RECT 5.635 0.265 5.92 0.965 ;
      RECT 6.495 0.265 6.825 0.855 ;
      RECT 5.635 0.265 6.825 0.435 ;
      RECT 6.115 2.015 6.445 2.735 ;
      RECT 5.4 2.015 6.445 2.205 ;
      RECT 1.355 2.905 3.19 3.075 ;
      RECT 3.02 2.035 3.19 3.075 ;
      RECT 2.295 1.03 2.465 3.075 ;
      RECT 1.355 2.63 1.615 3.075 ;
      RECT 5.605 2.375 5.935 2.735 ;
      RECT 3.02 2.375 5.935 2.545 ;
      RECT 3.02 2.035 3.69 2.545 ;
      RECT 3.52 0.295 3.69 2.545 ;
      RECT 4.37 1.335 6.325 1.505 ;
      RECT 6.09 0.645 6.325 1.505 ;
      RECT 4.37 0.295 4.54 1.505 ;
      RECT 0.975 1.03 2.465 1.215 ;
      RECT 0.885 0.645 1.215 1.03 ;
      RECT 3.52 0.295 4.54 0.465 ;
      RECT 2.635 0.58 2.85 2.735 ;
      RECT 2.295 0.58 2.85 0.86 ;
      RECT 0.095 2.29 0.425 3.075 ;
      RECT 1.785 2.29 2.115 2.735 ;
      RECT 0.095 2.29 2.115 2.46 ;
  END
END scs130lp_sdfxbp_2

MACRO scs130lp_sdfxbp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfxbp_lp 0 0 ;
  SIZE 15.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.485 1.18 4.195 1.51 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.925 1.215 2.275 1.885 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3963 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.125 1.985 12.835 3.025 ;
        RECT 12.125 1.125 12.76 1.295 ;
        RECT 12.51 0.615 12.76 1.295 ;
        RECT 12.125 1.125 12.295 3.025 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3984 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.715 1.92 15.74 3.065 ;
        RECT 15.41 0.265 15.74 3.065 ;
    END
  END QN
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.955 1.245 3.285 1.915 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.53 1.515 0.86 1.845 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 15.84 0.085 ;
        RECT 14.62 -0.085 14.95 0.725 ;
        RECT 13.3 -0.085 13.63 1.075 ;
        RECT 11.28 -0.085 11.53 0.595 ;
        RECT 7.85 -0.085 8.18 0.715 ;
        RECT 4.28 -0.085 4.61 0.65 ;
        RECT 2.95 -0.085 3.28 1.065 ;
        RECT 1.15 -0.085 1.48 0.985 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 15.84 3.415 ;
        RECT 14.185 2.335 14.515 3.415 ;
        RECT 13.015 1.985 13.345 3.415 ;
        RECT 10.75 2.13 11.08 3.415 ;
        RECT 7.875 2.015 8.205 3.415 ;
        RECT 4.32 2.505 4.65 3.415 ;
        RECT 2.69 2.855 3.02 3.415 ;
        RECT 0.63 2.025 0.96 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 13.545 1.985 13.875 3.025 ;
      RECT 13.545 1.985 14.515 2.155 ;
      RECT 14.345 0.905 14.515 2.155 ;
      RECT 14.345 0.905 14.825 1.575 ;
      RECT 14.09 0.615 14.42 1.075 ;
      RECT 11.36 2.13 11.69 2.825 ;
      RECT 11.36 2.13 11.9 2.3 ;
      RECT 11.73 0.775 11.9 2.3 ;
      RECT 12.475 1.475 14.165 1.805 ;
      RECT 10.565 0.965 10.895 1.6 ;
      RECT 12.94 0.265 13.11 1.805 ;
      RECT 10.565 0.965 11.9 1.135 ;
      RECT 11.73 0.775 12.32 0.945 ;
      RECT 11.99 0.265 12.32 0.945 ;
      RECT 11.99 0.265 13.11 0.435 ;
      RECT 9.565 1.715 9.895 2.78 ;
      RECT 9.565 1.78 11.55 1.95 ;
      RECT 11.22 1.315 11.55 1.95 ;
      RECT 9.75 0.965 10.08 1.95 ;
      RECT 9.255 0.615 9.505 1.215 ;
      RECT 9.255 0.615 11.1 0.785 ;
      RECT 10.77 0.265 11.1 0.785 ;
      RECT 8.745 0.265 9.075 2.755 ;
      RECT 7.65 1.155 7.98 1.485 ;
      RECT 7.81 0.895 7.98 1.485 ;
      RECT 7.81 0.895 9.075 1.065 ;
      RECT 8.705 0.265 9.075 1.065 ;
      RECT 8.705 0.265 10.575 0.435 ;
      RECT 6.855 1.395 7.185 2.755 ;
      RECT 6.855 1.665 8.55 1.835 ;
      RECT 8.22 1.245 8.55 1.835 ;
      RECT 6.375 1.395 7.185 1.565 ;
      RECT 6.375 0.965 6.705 1.565 ;
      RECT 5.595 0.265 5.845 1.125 ;
      RECT 7.355 0.265 7.605 0.975 ;
      RECT 5.595 0.265 7.605 0.435 ;
      RECT 6.025 1.745 6.655 2.755 ;
      RECT 1.69 2.155 6.655 2.325 ;
      RECT 1.69 2.065 2.625 2.325 ;
      RECT 2.455 0.605 2.625 2.325 ;
      RECT 6.025 0.615 6.195 2.755 ;
      RECT 6.885 0.615 7.135 1.215 ;
      RECT 2.16 0.605 2.625 1.035 ;
      RECT 6.025 0.615 7.135 0.785 ;
      RECT 4.85 1.715 5.66 1.975 ;
      RECT 5.23 1.305 5.66 1.975 ;
      RECT 5.23 0.31 5.4 1.975 ;
      RECT 5.07 0.31 5.4 0.65 ;
      RECT 3.79 1.715 4.545 1.975 ;
      RECT 4.375 0.83 4.545 1.975 ;
      RECT 4.375 0.83 4.91 1.53 ;
      RECT 3.49 0.83 4.91 1 ;
      RECT 3.49 0.31 3.82 1 ;
      RECT 3.22 2.505 3.55 3.065 ;
      RECT 1.16 2.065 1.49 3.065 ;
      RECT 1.16 2.505 3.55 2.675 ;
      RECT 0.1 0.605 0.35 3.065 ;
      RECT 1.355 1.165 1.685 1.835 ;
      RECT 0.1 1.165 1.685 1.335 ;
      RECT 0.1 0.605 0.58 1.335 ;
  END
END scs130lp_sdfxbp_lp

MACRO scs130lp_sdfxtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfxtp_1 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.255 1.175 3.695 2.215 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.455 0.385 1.775 2.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.195 0.365 10.465 3.075 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.985 1.495 2.735 1.795 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.445 1.145 1.285 1.475 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.56 0.085 ;
        RECT 9.74 -0.085 10.025 1.245 ;
        RECT 8.81 -0.085 9.02 0.975 ;
        RECT 6.225 -0.085 6.555 0.635 ;
        RECT 3.66 -0.085 3.92 0.545 ;
        RECT 2.655 -0.085 2.945 0.935 ;
        RECT 0.84 -0.085 1.05 0.925 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.56 3.415 ;
        RECT 9.74 1.815 9.975 3.415 ;
        RECT 8.755 2.345 9.085 3.415 ;
        RECT 6.33 2.975 6.66 3.415 ;
        RECT 3.635 2.725 3.895 3.415 ;
        RECT 2.755 2.66 2.945 3.415 ;
        RECT 0.95 2.64 1.245 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 4.895 2.29 5.185 2.52 ;
      RECT 2.495 2.29 2.785 2.52 ;
      RECT 2.495 2.335 5.185 2.475 ;
    LAYER li ;
      RECT 9.265 1.985 9.57 2.91 ;
      RECT 9.4 0.315 9.57 2.91 ;
      RECT 8.285 1.985 9.57 2.175 ;
      RECT 9.4 1.415 9.78 1.645 ;
      RECT 9.24 0.315 9.57 0.985 ;
      RECT 7.69 2.515 7.955 2.845 ;
      RECT 7.785 1.645 7.955 2.845 ;
      RECT 7.785 1.645 9.22 1.815 ;
      RECT 8.42 1.305 9.22 1.815 ;
      RECT 8.42 0.345 8.59 1.815 ;
      RECT 7.945 0.345 8.59 0.675 ;
      RECT 4.065 2.895 5.93 3.065 ;
      RECT 5.76 1.515 5.93 3.065 ;
      RECT 3.115 2.385 3.445 3.045 ;
      RECT 4.065 0.715 4.235 3.065 ;
      RECT 5.76 2.635 7.52 2.805 ;
      RECT 7.35 1.755 7.52 2.805 ;
      RECT 3.115 2.385 4.235 2.555 ;
      RECT 3.865 0.715 4.235 2.555 ;
      RECT 7.435 1.295 7.605 2.085 ;
      RECT 5.465 1.515 5.93 1.705 ;
      RECT 7.435 1.295 8.25 1.465 ;
      RECT 7.99 0.855 8.25 1.465 ;
      RECT 3.115 0.715 4.235 0.985 ;
      RECT 4.405 0.265 4.595 2.725 ;
      RECT 7.435 0.385 7.765 1.125 ;
      RECT 5.68 0.815 6.905 0.985 ;
      RECT 6.735 0.385 6.905 0.985 ;
      RECT 5.68 0.265 5.85 0.985 ;
      RECT 6.735 0.385 7.765 0.555 ;
      RECT 4.09 0.265 5.85 0.485 ;
      RECT 6.1 1.685 7.17 2.465 ;
      RECT 7 1.165 7.17 2.465 ;
      RECT 7.075 0.735 7.265 1.335 ;
      RECT 5.34 1.875 5.59 2.615 ;
      RECT 5.115 1.875 5.59 2.045 ;
      RECT 5.115 1.175 5.285 2.045 ;
      RECT 6.65 1.175 6.82 1.505 ;
      RECT 5.115 1.175 6.82 1.345 ;
      RECT 5.265 0.655 5.51 1.345 ;
      RECT 4.765 2.225 5.17 2.555 ;
      RECT 4.765 0.665 4.935 2.555 ;
      RECT 4.765 0.665 5.095 0.995 ;
      RECT 1.75 2.64 2.585 2.97 ;
      RECT 2.415 2.035 2.585 2.97 ;
      RECT 2.415 2.035 2.725 2.49 ;
      RECT 2.415 2.035 3.075 2.205 ;
      RECT 2.905 1.155 3.075 2.205 ;
      RECT 1.945 1.155 3.075 1.325 ;
      RECT 1.945 0.685 2.195 1.325 ;
      RECT 0.45 1.655 0.78 3.045 ;
      RECT 0.45 2.3 2.235 2.47 ;
      RECT 1.995 1.965 2.235 2.47 ;
      RECT 0.45 1.655 1.235 2.47 ;
      RECT 0.095 1.655 1.235 1.985 ;
      RECT 0.095 0.635 0.265 1.985 ;
      RECT 0.095 0.635 0.62 0.965 ;
  END
END scs130lp_sdfxtp_1

MACRO scs130lp_sdfxtp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfxtp_2 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.255 1.2 3.735 2.12 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.115 0.385 1.765 1.455 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.225 0.375 10.465 3.075 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.035 1.455 2.725 1.775 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.45 1.14 0.83 2.13 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 10.635 -0.085 10.935 1.255 ;
        RECT 9.745 -0.085 10.055 1.175 ;
        RECT 8.83 -0.085 9.04 0.885 ;
        RECT 6.205 -0.085 6.545 0.555 ;
        RECT 3.695 -0.085 4.025 0.53 ;
        RECT 2.695 -0.085 3.025 0.945 ;
        RECT 0.725 -0.085 0.945 0.97 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.04 3.415 ;
        RECT 10.635 1.815 10.935 3.415 ;
        RECT 9.745 1.845 10.055 3.415 ;
        RECT 8.45 2.325 9.125 3.415 ;
        RECT 6.095 2.455 6.375 3.415 ;
        RECT 3.555 2.64 3.805 3.415 ;
        RECT 2.625 2.69 2.845 3.415 ;
        RECT 0.78 2.64 1.11 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 4.895 2.29 5.185 2.52 ;
      RECT 2.495 2.29 2.785 2.52 ;
      RECT 2.495 2.335 5.185 2.475 ;
    LAYER li ;
      RECT 9.295 1.975 9.55 2.905 ;
      RECT 9.38 0.255 9.55 2.905 ;
      RECT 8.325 1.975 9.55 2.155 ;
      RECT 9.38 1.345 10.055 1.675 ;
      RECT 9.21 0.255 9.55 0.895 ;
      RECT 7.635 2.235 7.985 3.075 ;
      RECT 7.815 1.635 7.985 3.075 ;
      RECT 7.815 1.635 9.21 1.805 ;
      RECT 8.49 1.135 9.21 1.805 ;
      RECT 8.49 0.335 8.66 1.805 ;
      RECT 7.975 0.335 8.66 0.665 ;
      RECT 3.025 2.3 3.355 3.025 ;
      RECT 3.975 2.835 5.845 3.005 ;
      RECT 5.675 1.425 5.845 3.005 ;
      RECT 6.545 2.745 7.465 2.915 ;
      RECT 3.975 0.86 4.145 3.005 ;
      RECT 7.295 1.835 7.465 2.915 ;
      RECT 6.545 2.115 6.715 2.915 ;
      RECT 3.025 2.3 4.145 2.47 ;
      RECT 3.905 0.86 4.145 2.47 ;
      RECT 5.675 2.115 6.715 2.285 ;
      RECT 7.465 1.275 7.635 2.065 ;
      RECT 5.485 1.425 5.845 1.755 ;
      RECT 7.465 1.275 8.32 1.445 ;
      RECT 8.02 0.845 8.32 1.445 ;
      RECT 3.225 0.7 3.905 1.03 ;
      RECT 4.315 1.175 4.625 2.665 ;
      RECT 4.315 0.265 4.535 2.665 ;
      RECT 7.465 0.255 7.795 1.095 ;
      RECT 5.66 0.725 6.935 0.895 ;
      RECT 6.715 0.255 6.935 0.895 ;
      RECT 5.66 0.265 5.965 0.895 ;
      RECT 4.195 0.265 4.535 0.61 ;
      RECT 4.195 0.265 5.965 0.485 ;
      RECT 6.715 0.255 7.795 0.425 ;
      RECT 6.885 1.495 7.125 2.575 ;
      RECT 6.025 1.495 7.125 1.945 ;
      RECT 7.105 0.595 7.295 1.665 ;
      RECT 6.025 1.425 6.355 1.945 ;
      RECT 5.305 1.935 5.495 2.63 ;
      RECT 5.145 1.075 5.315 2.105 ;
      RECT 6.605 1.075 6.935 1.325 ;
      RECT 5.145 1.075 6.935 1.245 ;
      RECT 5.27 0.67 5.49 1.245 ;
      RECT 4.795 2.275 5.135 2.59 ;
      RECT 4.795 0.655 4.965 2.59 ;
      RECT 4.76 0.655 4.965 0.955 ;
      RECT 4.76 0.655 5.09 0.905 ;
      RECT 1.615 2.445 1.945 3.075 ;
      RECT 1.615 2.445 2.455 2.645 ;
      RECT 2.285 1.95 2.725 2.52 ;
      RECT 2.285 1.95 3.075 2.12 ;
      RECT 2.905 1.115 3.075 2.12 ;
      RECT 1.935 1.115 3.075 1.285 ;
      RECT 1.935 0.635 2.135 1.285 ;
      RECT 0.315 2.3 0.61 3.075 ;
      RECT 0.11 2.3 1.17 2.47 ;
      RECT 1 1.635 1.17 2.47 ;
      RECT 0.11 0.64 0.28 2.47 ;
      RECT 1 1.945 2.115 2.275 ;
      RECT 1 1.635 1.25 2.275 ;
      RECT 0.11 0.64 0.555 0.97 ;
  END
END scs130lp_sdfxtp_2

MACRO scs130lp_sdfxtp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfxtp_4 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.255 1.19 3.695 2.12 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.51 0.47 1.775 2.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.205 0.945 11.91 1.925 ;
        RECT 11.205 0.255 11.395 3.075 ;
        RECT 10.31 1.655 11.91 1.825 ;
        RECT 11.195 0.945 11.91 1.825 ;
        RECT 10.305 0.945 11.91 1.115 ;
        RECT 10.31 1.655 10.535 3.075 ;
        RECT 10.305 0.255 10.535 1.115 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.945 1.395 2.725 1.795 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.48 1.145 1.34 1.475 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12 0.085 ;
        RECT 11.565 -0.085 11.895 0.775 ;
        RECT 10.705 -0.085 11.035 0.775 ;
        RECT 9.845 -0.085 10.135 1.115 ;
        RECT 8.855 -0.085 9.175 1.015 ;
        RECT 6.255 -0.085 6.585 0.385 ;
        RECT 3.795 -0.085 4.125 0.615 ;
        RECT 2.75 -0.085 3.08 0.875 ;
        RECT 0.845 -0.085 1.175 0.975 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
      LAYER li ;
        RECT 0 3.245 12 3.415 ;
        RECT 11.565 2.095 11.895 3.415 ;
        RECT 10.705 1.995 11.035 3.415 ;
        RECT 9.845 1.815 10.14 3.415 ;
        RECT 8.495 2.58 9.225 3.415 ;
        RECT 8.895 2.405 9.225 3.415 ;
        RECT 6.41 2.975 6.74 3.415 ;
        RECT 3.7 2.64 3.96 3.415 ;
        RECT 2.82 2.66 3.01 3.415 ;
        RECT 1.025 2.64 1.355 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 4.895 2.29 5.185 2.52 ;
      RECT 2.495 2.29 2.785 2.52 ;
      RECT 2.495 2.335 5.185 2.475 ;
    LAYER li ;
      RECT 9.395 2.045 9.595 2.975 ;
      RECT 9.405 0.255 9.595 2.975 ;
      RECT 8.495 2.045 8.725 2.375 ;
      RECT 8.495 2.045 9.595 2.215 ;
      RECT 9.405 1.285 11.015 1.485 ;
      RECT 9.405 0.255 9.605 1.485 ;
      RECT 9.345 0.255 9.605 1.005 ;
      RECT 7.77 2.58 8.325 2.91 ;
      RECT 8.155 1.695 8.325 2.91 ;
      RECT 8.155 1.695 8.685 1.865 ;
      RECT 8.515 0.345 8.685 1.865 ;
      RECT 8.515 1.185 9.235 1.515 ;
      RECT 7.965 0.345 8.685 0.675 ;
      RECT 3.18 2.505 3.51 3.075 ;
      RECT 3.34 2.3 3.51 3.075 ;
      RECT 4.13 2.895 6.045 3.065 ;
      RECT 5.875 1.515 6.045 3.065 ;
      RECT 4.13 0.785 4.3 3.065 ;
      RECT 5.875 2.635 7.6 2.805 ;
      RECT 7.43 1.825 7.6 2.805 ;
      RECT 3.34 2.3 4.3 2.47 ;
      RECT 3.865 0.785 4.3 2.47 ;
      RECT 7.27 1.825 7.6 2.035 ;
      RECT 7.27 1.825 7.975 2.005 ;
      RECT 5.71 1.515 6.045 1.845 ;
      RECT 7.805 1.345 7.975 2.005 ;
      RECT 7.975 0.855 8.335 1.515 ;
      RECT 3.275 0.785 4.3 1.02 ;
      RECT 4.47 1.235 4.75 2.725 ;
      RECT 4.47 0.255 4.665 2.725 ;
      RECT 7.615 0.255 7.795 1.165 ;
      RECT 5.72 0.555 6.935 0.725 ;
      RECT 6.765 0.255 6.935 0.725 ;
      RECT 4.295 0.255 4.665 0.595 ;
      RECT 5.72 0.255 5.89 0.725 ;
      RECT 4.295 0.255 5.89 0.495 ;
      RECT 6.765 0.255 7.795 0.425 ;
      RECT 6.92 2.205 7.25 2.465 ;
      RECT 6.92 1.475 7.09 2.465 ;
      RECT 6.225 1.475 7.09 2.075 ;
      RECT 6.225 1.475 7.445 1.655 ;
      RECT 7.275 0.595 7.445 1.655 ;
      RECT 7.115 0.595 7.445 0.885 ;
      RECT 5.36 2.225 5.705 2.725 ;
      RECT 5.36 0.665 5.54 2.725 ;
      RECT 5.36 1.055 7.095 1.305 ;
      RECT 5.32 0.665 5.55 1.12 ;
      RECT 4.92 2.295 5.19 2.625 ;
      RECT 4.92 0.665 5.15 2.625 ;
      RECT 4.835 0.665 5.15 0.995 ;
      RECT 1.815 2.64 2.65 2.97 ;
      RECT 2.48 2.155 2.65 2.97 ;
      RECT 2.48 2.155 3.01 2.49 ;
      RECT 2.905 1.045 3.075 2.335 ;
      RECT 1.945 1.045 3.075 1.215 ;
      RECT 1.945 0.725 2.135 1.215 ;
      RECT 0.13 1.655 0.855 2.945 ;
      RECT 0.13 2.3 2.31 2.47 ;
      RECT 2.05 1.965 2.31 2.47 ;
      RECT 0.13 1.655 1.27 2.47 ;
      RECT 0.13 0.635 0.31 2.945 ;
      RECT 0.13 0.635 0.675 0.965 ;
  END
END scs130lp_sdfxtp_4

MACRO scs130lp_sdfxtp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdfxtp_lp 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.95 1.18 4.28 1.51 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.965 1.215 2.295 1.885 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.605 1.92 13.275 2.96 ;
        RECT 12.905 0.325 13.075 2.96 ;
        RECT 12.685 0.325 13.075 0.785 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.313 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.005 1.245 3.715 1.915 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 1.515 0.875 1.845 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.92 0.085 ;
        RECT 13.475 -0.085 13.805 0.785 ;
        RECT 11.34 -0.085 11.67 0.785 ;
        RECT 8.08 -0.085 8.41 0.715 ;
        RECT 4.435 -0.085 4.765 0.65 ;
        RECT 3.09 -0.085 3.42 1.065 ;
        RECT 1.16 -0.085 1.49 0.985 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.92 3.415 ;
        RECT 13.475 1.92 13.805 3.415 ;
        RECT 10.965 1.825 11.295 3.415 ;
        RECT 8.105 2.015 8.435 3.415 ;
        RECT 4.435 2.505 4.765 3.415 ;
        RECT 2.73 2.855 3.06 3.415 ;
        RECT 0.645 2.025 0.975 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 11.57 1.825 12.025 2.825 ;
      RECT 11.855 0.965 12.025 2.825 ;
      RECT 12.395 0.965 12.725 1.635 ;
      RECT 10.775 0.965 11.105 1.295 ;
      RECT 10.775 0.965 12.725 1.135 ;
      RECT 12.13 0.325 12.3 1.135 ;
      RECT 12.13 0.325 12.46 0.785 ;
      RECT 9.84 1.475 10.17 2.825 ;
      RECT 9.84 1.475 11.675 1.645 ;
      RECT 11.345 1.315 11.675 1.645 ;
      RECT 9.94 0.965 10.27 1.645 ;
      RECT 9.53 0.615 9.77 1.215 ;
      RECT 9.53 0.615 11.16 0.785 ;
      RECT 10.91 0.325 11.16 0.785 ;
      RECT 9.105 1.715 9.435 2.755 ;
      RECT 9.105 0.265 9.275 2.755 ;
      RECT 7.88 1.155 8.21 1.485 ;
      RECT 8.04 0.895 8.21 1.485 ;
      RECT 8.04 0.895 9.275 1.065 ;
      RECT 8.945 0.265 9.275 1.065 ;
      RECT 8.945 0.265 10.685 0.435 ;
      RECT 7.085 1.365 7.415 2.755 ;
      RECT 7.085 1.665 8.79 1.835 ;
      RECT 8.46 1.245 8.79 1.835 ;
      RECT 6.56 1.365 7.415 1.535 ;
      RECT 6.56 0.965 6.89 1.535 ;
      RECT 5.78 0.265 6.03 1.125 ;
      RECT 7.575 0.265 7.825 0.975 ;
      RECT 5.78 0.265 7.825 0.435 ;
      RECT 6.555 1.715 6.885 2.755 ;
      RECT 1.73 2.155 6.885 2.325 ;
      RECT 6.21 1.715 6.885 2.325 ;
      RECT 1.73 2.065 2.645 2.325 ;
      RECT 2.475 0.605 2.645 2.325 ;
      RECT 6.21 0.615 6.38 2.325 ;
      RECT 7.07 0.615 7.32 1.185 ;
      RECT 2.2 0.605 2.645 1.035 ;
      RECT 6.21 0.615 7.32 0.785 ;
      RECT 4.965 1.715 5.82 1.975 ;
      RECT 5.225 1.305 5.82 1.975 ;
      RECT 5.225 0.31 5.555 1.975 ;
      RECT 3.905 1.715 4.63 1.975 ;
      RECT 4.46 0.83 4.63 1.975 ;
      RECT 4.46 0.83 5.045 1.53 ;
      RECT 3.645 0.83 5.045 1 ;
      RECT 3.645 0.31 3.975 1 ;
      RECT 3.26 2.505 3.59 3.065 ;
      RECT 1.2 2.065 1.53 3.065 ;
      RECT 1.2 2.505 3.59 2.675 ;
      RECT 0.115 0.605 0.365 3.065 ;
      RECT 1.425 1.165 1.755 1.835 ;
      RECT 0.115 1.165 1.755 1.335 ;
      RECT 0.115 0.605 0.67 1.335 ;
  END
END scs130lp_sdfxtp_lp

MACRO scs130lp_sdlclkp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdlclkp_1 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.64 0.805 6.195 1.39 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.06 0.84 1.365 1.76 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 0.5565 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.15 1.85 7.595 3.075 ;
        RECT 7.325 0.255 7.595 3.075 ;
    END
  END GCLK
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.465 2.49 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
      LAYER li ;
        RECT 0 -0.085 7.68 0.085 ;
        RECT 6.825 -0.085 7.155 0.815 ;
        RECT 5.575 -0.085 5.785 0.635 ;
        RECT 4.02 -0.085 4.35 0.355 ;
        RECT 1.245 -0.085 1.475 0.67 ;
        RECT 0.29 -0.085 0.54 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
      LAYER li ;
        RECT 0 3.245 7.68 3.415 ;
        RECT 6.64 2.25 6.97 3.415 ;
        RECT 5.62 2.565 5.95 3.415 ;
        RECT 4.135 1.985 4.465 3.415 ;
        RECT 1.455 2.27 1.715 3.415 ;
        RECT 0.095 2.66 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.13 1.91 6.46 2.44 ;
      RECT 6.13 1.91 6.97 2.08 ;
      RECT 6.8 0.985 6.97 2.08 ;
      RECT 6.8 1.185 7.155 1.515 ;
      RECT 6.365 0.985 6.97 1.155 ;
      RECT 6.365 0.305 6.635 1.155 ;
      RECT 4.635 1.645 4.93 3.075 ;
      RECT 4.76 0.865 4.93 3.075 ;
      RECT 4.635 2.225 5.79 2.395 ;
      RECT 5.62 1.56 5.79 2.395 ;
      RECT 3.685 1.645 3.965 1.975 ;
      RECT 3.685 1.645 4.93 1.815 ;
      RECT 5.62 1.56 6.63 1.73 ;
      RECT 6.365 1.345 6.63 1.73 ;
      RECT 4.53 0.865 4.93 1.105 ;
      RECT 5.11 1.795 5.44 2.055 ;
      RECT 5.11 0.305 5.355 2.055 ;
      RECT 2.145 0.37 2.405 1.345 ;
      RECT 3.68 0.525 5.355 0.695 ;
      RECT 5.085 0.305 5.355 0.695 ;
      RECT 2.145 0.37 3.85 0.54 ;
      RECT 3.255 0.71 3.495 2.69 ;
      RECT 3.255 1.275 4.58 1.475 ;
      RECT 3.14 0.71 3.495 1.33 ;
      RECT 1.885 2.875 3.085 3.045 ;
      RECT 2.8 1.5 3.085 3.045 ;
      RECT 0.71 1.93 1.215 2.99 ;
      RECT 1.885 1.93 2.055 3.045 ;
      RECT 0.71 1.93 2.055 2.1 ;
      RECT 0.71 0.39 0.88 2.99 ;
      RECT 2.8 0.71 2.97 3.045 ;
      RECT 2.64 0.71 2.97 1.04 ;
      RECT 0.71 0.39 1.075 0.67 ;
      RECT 2.225 1.555 2.475 2.695 ;
      RECT 2.225 1.555 2.63 1.885 ;
      RECT 1.645 1.555 2.63 1.76 ;
      RECT 1.645 0.39 1.975 1.76 ;
  END
END scs130lp_sdlclkp_1

MACRO scs130lp_sdlclkp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdlclkp_2 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.415 0.84 5.79 1.565 ;
        RECT 5.415 0.84 5.615 1.83 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.925 1.305 1.315 1.975 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 0.588 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.285 1.855 7.615 2.045 ;
        RECT 7.345 0.255 7.615 2.045 ;
    END
  END GCLK
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.415 2.16 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.785 -0.085 8.045 1.125 ;
        RECT 6.845 -0.085 7.175 0.875 ;
        RECT 5.415 -0.085 5.745 0.67 ;
        RECT 3.915 -0.085 4.245 0.355 ;
        RECT 0.99 -0.085 1.25 0.725 ;
        RECT 0.095 -0.085 0.425 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.715 2.555 8.045 3.415 ;
        RECT 6.58 2.555 7.185 3.415 ;
        RECT 5.64 2.875 5.97 3.415 ;
        RECT 4.045 2.085 4.49 3.415 ;
        RECT 1.465 2.505 1.795 3.415 ;
        RECT 0.095 2.33 0.415 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.15 2.075 6.41 2.825 ;
      RECT 6.15 2.215 8.045 2.385 ;
      RECT 7.785 1.295 8.045 2.385 ;
      RECT 6.15 2.075 7.115 2.385 ;
      RECT 6.895 1.045 7.115 2.385 ;
      RECT 6.205 1.045 7.115 1.215 ;
      RECT 6.205 0.45 6.535 1.215 ;
      RECT 4.66 2.535 4.92 3.075 ;
      RECT 4.66 2.535 5.955 2.705 ;
      RECT 5.785 1.735 5.955 2.705 ;
      RECT 4.66 1.745 4.9 3.075 ;
      RECT 4.73 0.865 4.9 3.075 ;
      RECT 3.715 1.745 4.9 1.915 ;
      RECT 5.785 1.735 6.715 1.905 ;
      RECT 6.385 1.385 6.715 1.905 ;
      RECT 3.715 1.585 4.04 1.915 ;
      RECT 4.425 0.865 4.9 1.055 ;
      RECT 5.07 2.115 5.46 2.365 ;
      RECT 5.07 0.365 5.245 2.365 ;
      RECT 1.905 0.255 2.235 0.855 ;
      RECT 1.905 0.525 5.245 0.695 ;
      RECT 4.985 0.365 5.245 0.695 ;
      RECT 3.305 0.865 3.545 2.655 ;
      RECT 4.3 1.225 4.56 1.555 ;
      RECT 3.045 1.225 4.56 1.395 ;
      RECT 3.045 0.865 3.545 1.395 ;
      RECT 1.965 2.895 3.135 3.065 ;
      RECT 2.695 2.325 3.135 3.065 ;
      RECT 0.585 2.165 1.215 2.99 ;
      RECT 1.965 2.165 2.135 3.065 ;
      RECT 0.585 2.165 2.135 2.335 ;
      RECT 2.695 0.865 2.865 3.065 ;
      RECT 0.585 0.74 0.755 2.99 ;
      RECT 2.535 0.865 2.865 1.125 ;
      RECT 0.595 0.395 0.82 0.93 ;
      RECT 2.305 1.585 2.525 2.725 ;
      RECT 1.485 1.585 2.525 1.915 ;
      RECT 1.485 0.395 1.715 1.915 ;
      RECT 1.42 0.395 1.715 1.125 ;
  END
END scs130lp_sdlclkp_2

MACRO scs130lp_sdlclkp_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdlclkp_4 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.474 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.435 1.21 6.085 1.76 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.065 1.045 2.245 1.79 ;
        RECT 1.065 0.925 1.315 1.79 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 1.176 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.305 0.425 8.505 2.47 ;
        RECT 8.21 1.605 8.445 3.075 ;
        RECT 7.445 0.845 8.505 1.015 ;
        RECT 7.365 1.605 8.505 1.775 ;
        RECT 7.445 0.255 7.635 1.015 ;
        RECT 7.365 1.605 7.61 3.075 ;
    END
  END GCLK
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 0.84 0.435 2.49 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 8.675 -0.085 8.995 1.09 ;
        RECT 7.805 -0.085 8.135 0.675 ;
        RECT 6.945 -0.085 7.275 0.825 ;
        RECT 5.625 -0.085 5.955 1.04 ;
        RECT 4.05 -0.085 4.38 0.355 ;
        RECT 1.17 -0.085 1.48 0.725 ;
        RECT 0.205 -0.085 0.535 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 8.675 1.815 8.935 3.415 ;
        RECT 7.78 1.945 8.04 3.415 ;
        RECT 6.955 2.185 7.195 3.415 ;
        RECT 5.98 2.785 6.19 3.415 ;
        RECT 3.935 2.36 4.53 3.415 ;
        RECT 4.34 1.985 4.53 3.415 ;
        RECT 1.445 2.3 1.705 3.415 ;
        RECT 0.095 2.66 0.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.41 2.28 6.785 2.95 ;
      RECT 6.615 1.845 6.785 2.95 ;
      RECT 6.615 1.845 7.195 2.015 ;
      RECT 7.025 0.995 7.195 2.015 ;
      RECT 7.025 1.185 8.135 1.435 ;
      RECT 6.415 0.995 7.195 1.175 ;
      RECT 6.415 0.255 6.685 1.175 ;
      RECT 4.71 2.31 5.04 2.93 ;
      RECT 4.71 2.31 6.075 2.49 ;
      RECT 5.905 1.93 6.075 2.49 ;
      RECT 4.71 1.635 4.915 2.93 ;
      RECT 4.72 0.865 4.915 2.93 ;
      RECT 5.905 1.93 6.435 2.1 ;
      RECT 6.265 1.345 6.435 2.1 ;
      RECT 3.805 1.635 4.14 2.095 ;
      RECT 3.805 1.635 4.915 1.805 ;
      RECT 6.265 1.345 6.855 1.675 ;
      RECT 4.56 0.865 4.915 1.08 ;
      RECT 5.085 1.93 5.725 2.14 ;
      RECT 5.085 0.27 5.255 2.14 ;
      RECT 3.7 0.525 5.43 0.695 ;
      RECT 5.085 0.27 5.43 0.695 ;
      RECT 3.7 0.255 3.87 0.695 ;
      RECT 2.265 0.255 3.87 0.445 ;
      RECT 3.18 0.71 3.475 2.695 ;
      RECT 3.18 1.25 4.54 1.465 ;
      RECT 1.875 2.885 3.01 3.075 ;
      RECT 2.775 0.71 3.01 3.075 ;
      RECT 0.705 1.96 1.215 2.99 ;
      RECT 1.875 1.96 2.045 3.075 ;
      RECT 0.705 1.96 2.045 2.13 ;
      RECT 0.705 0.395 0.895 2.99 ;
      RECT 0.705 0.395 0.975 0.725 ;
      RECT 2.225 2.045 2.605 2.715 ;
      RECT 2.425 0.615 2.605 2.715 ;
      RECT 1.65 0.615 2.605 0.785 ;
      RECT 1.65 0.395 1.98 0.785 ;
  END
END scs130lp_sdlclkp_4

MACRO scs130lp_sdlclkp_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sdlclkp_lp 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 4.925 1.58 5.655 2.15 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.035 0.555 1.705 ;
    END
  END GATE
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.115 2.06 8.515 3.065 ;
        RECT 8.285 0.265 8.515 3.065 ;
        RECT 8.075 0.265 8.515 0.595 ;
    END
  END GCLK
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.39 1.57 2.15 ;
    END
  END SCE
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.64 0.085 ;
        RECT 7.265 -0.085 7.595 0.68 ;
        RECT 6.585 -0.085 6.835 1.4 ;
        RECT 4.425 -0.085 4.755 0.675 ;
        RECT 1.725 -0.085 2.055 0.86 ;
        RECT 0.115 -0.085 0.445 0.855 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.64 3.415 ;
        RECT 7.505 2.84 7.835 3.415 ;
        RECT 6.365 2.84 6.695 3.415 ;
        RECT 4.525 2.68 4.855 3.415 ;
        RECT 1.545 2.965 1.875 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.895 2.06 7.225 2.31 ;
      RECT 6.895 2.06 7.575 2.23 ;
      RECT 7.325 0.935 7.575 2.23 ;
      RECT 7.325 0.935 8.105 1.105 ;
      RECT 7.775 0.775 8.105 1.105 ;
      RECT 5.09 2.33 5.42 3.045 ;
      RECT 5.09 2.49 7.925 2.66 ;
      RECT 7.755 1.315 7.925 2.66 ;
      RECT 4.325 2.33 5.42 2.5 ;
      RECT 6.345 1.58 6.515 2.66 ;
      RECT 4.325 1.58 4.655 2.5 ;
      RECT 6.225 0.505 6.395 1.75 ;
      RECT 7.755 1.315 8.085 1.645 ;
      RECT 5.445 0.505 6.395 0.675 ;
      RECT 5.445 0.265 5.775 0.675 ;
      RECT 2.405 2.435 4.145 2.605 ;
      RECT 3.975 1.23 4.145 2.605 ;
      RECT 1.78 2.265 2.575 2.435 ;
      RECT 5.835 2.06 6.165 2.31 ;
      RECT 1.78 1.39 2.11 2.435 ;
      RECT 5.835 0.94 6.045 2.31 ;
      RECT 3.73 1.495 4.145 1.825 ;
      RECT 3.975 1.23 6.045 1.4 ;
      RECT 5.715 0.94 6.045 1.4 ;
      RECT 3.38 2.005 3.795 2.255 ;
      RECT 3.38 0.88 3.55 2.255 ;
      RECT 3.38 0.88 5.265 1.05 ;
      RECT 4.935 0.765 5.265 1.05 ;
      RECT 3.685 0.265 3.935 1.05 ;
      RECT 2.055 2.785 3.265 3.045 ;
      RECT 0.445 1.885 0.775 2.9 ;
      RECT 0.445 2.615 2.225 2.785 ;
      RECT 0.735 0.485 0.905 2.785 ;
      RECT 0.735 1.04 2.405 1.21 ;
      RECT 2.235 0.265 2.405 1.21 ;
      RECT 0.735 0.485 1.265 1.21 ;
      RECT 3.175 0.265 3.505 0.675 ;
      RECT 2.235 0.265 3.505 0.435 ;
      RECT 2.29 1.39 2.62 2.085 ;
      RECT 2.29 1.39 3.2 1.72 ;
      RECT 2.8 0.615 2.97 1.72 ;
      RECT 2.595 0.615 2.97 0.945 ;
  END
END scs130lp_sdlclkp_lp

MACRO scs130lp_sleep_pargate_plv_14
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sleep_pargate_plv_14 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.1 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.8 8.785 2.83 ;
    END
  END sleep
  PIN virtpwr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855 LAYER li ;
    ANTENNADIFFAREA 3.71 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
        RECT 6.51 1.965 7.155 3.575 ;
        RECT 4.955 1.965 5.58 3.575 ;
        RECT 3.4 1.965 4.025 3.575 ;
        RECT 1.845 1.965 2.47 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 1.055 2.84 8.055 3.415 ;
        RECT 1.055 1.98 7.95 2.24 ;
    END
  END virtpwr
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.28 0 8.84 3.33 ;
      LAYER met1 ;
        RECT 7.295 2.41 7.945 2.67 ;
        RECT 5.72 2.41 6.37 2.67 ;
        RECT 4.165 2.41 4.815 2.67 ;
        RECT 2.61 2.41 3.26 2.67 ;
        RECT 1.055 2.41 1.705 2.67 ;
      LAYER li ;
        RECT 1.055 2.41 7.95 2.67 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
END scs130lp_sleep_pargate_plv_14

MACRO scs130lp_sleep_pargate_plv_21
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sleep_pargate_plv_21 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 3.15 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.8 8.785 2.83 ;
    END
  END sleep
  PIN virtpwr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855 LAYER li ;
    ANTENNADIFFAREA 3.815 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
        RECT 6.51 1.55 7.155 3.575 ;
        RECT 4.955 1.55 5.58 3.575 ;
        RECT 3.4 1.55 4.025 3.575 ;
        RECT 1.845 1.55 2.47 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 1.055 2.84 8.055 3.415 ;
        RECT 1.055 1.98 7.95 2.24 ;
    END
  END virtpwr
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.28 0 8.84 3.33 ;
      LAYER met1 ;
        RECT 7.295 1.55 7.945 2.67 ;
        RECT 5.72 1.55 6.37 2.67 ;
        RECT 4.165 1.55 4.815 2.67 ;
        RECT 2.61 1.55 3.26 2.67 ;
        RECT 1.055 1.55 1.705 2.67 ;
      LAYER li ;
        RECT 1.055 1.55 7.95 1.81 ;
        RECT 1.055 2.41 7.95 2.67 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
END scs130lp_sleep_pargate_plv_21

MACRO scs130lp_sleep_pargate_plv_28
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sleep_pargate_plv_28 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 4.2 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.8 8.785 2.83 ;
    END
  END sleep
  PIN virtpwr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855 LAYER li ;
    ANTENNADIFFAREA 5.95 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
        RECT 6.51 1.105 7.155 3.575 ;
        RECT 4.955 1.105 5.58 3.575 ;
        RECT 3.4 1.105 4.025 3.575 ;
        RECT 1.845 1.105 2.47 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 1.055 2.84 8.055 3.415 ;
        RECT 1.055 1.12 7.95 1.38 ;
        RECT 1.055 1.98 7.95 2.24 ;
    END
  END virtpwr
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.28 0 8.84 3.33 ;
      LAYER met1 ;
        RECT 7.295 1.55 7.945 2.67 ;
        RECT 5.72 1.55 6.37 2.67 ;
        RECT 4.165 1.55 4.815 2.67 ;
        RECT 2.61 1.55 3.26 2.67 ;
        RECT 1.055 1.55 1.705 2.67 ;
      LAYER li ;
        RECT 1.055 1.55 7.95 1.81 ;
        RECT 1.055 2.41 7.95 2.67 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
END scs130lp_sleep_pargate_plv_28

MACRO scs130lp_sleep_pargate_plv_7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sleep_pargate_plv_7 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.05 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.8 8.785 2.83 ;
    END
  END sleep
  PIN virtpwr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855 LAYER li ;
    ANTENNADIFFAREA 1.855 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
        RECT 6.51 2.825 7.155 3.575 ;
        RECT 4.955 2.825 5.58 3.575 ;
        RECT 3.4 2.825 4.025 3.575 ;
        RECT 1.845 2.825 2.47 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 1.055 2.84 8.055 3.415 ;
    END
  END virtpwr
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.28 0 8.84 3.33 ;
      LAYER met1 ;
        RECT 7.295 2.41 7.945 2.67 ;
        RECT 5.72 2.41 6.37 2.67 ;
        RECT 4.165 2.41 4.815 2.67 ;
        RECT 2.61 2.41 3.26 2.67 ;
        RECT 1.055 2.41 1.705 2.67 ;
      LAYER li ;
        RECT 1.055 2.41 7.95 2.67 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
END scs130lp_sleep_pargate_plv_7

MACRO scs130lp_sleep_sergate_plv_14
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sleep_sergate_plv_14 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.1 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.8 8.785 2.83 ;
    END
  END sleep
  PIN virtpwr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855 LAYER li ;
    ANTENNADIFFAREA 3.71 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
        RECT 6.51 1.965 7.155 3.575 ;
        RECT 4.955 1.965 5.58 3.575 ;
        RECT 3.4 1.965 4.025 3.575 ;
        RECT 1.845 1.965 2.47 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 1.055 2.84 8.055 3.415 ;
        RECT 1.055 1.98 7.95 2.24 ;
    END
  END virtpwr
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.295 2.41 7.945 2.67 ;
        RECT 5.72 2.41 6.37 2.67 ;
        RECT 4.165 2.41 4.815 2.67 ;
        RECT 2.61 2.41 3.26 2.67 ;
        RECT 1.055 2.41 1.705 2.67 ;
      LAYER met2 ;
        RECT 0.28 0 8.84 3.33 ;
      LAYER li ;
        RECT 1.055 2.41 7.95 2.67 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
END scs130lp_sleep_sergate_plv_14

MACRO scs130lp_sleep_sergate_plv_21
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sleep_sergate_plv_21 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 3.15 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.8 8.785 2.83 ;
    END
  END sleep
  PIN virtpwr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855 LAYER li ;
    ANTENNADIFFAREA 3.815 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
        RECT 6.51 1.55 7.155 3.575 ;
        RECT 4.955 1.55 5.58 3.575 ;
        RECT 3.4 1.55 4.025 3.575 ;
        RECT 1.845 1.55 2.47 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 1.055 2.84 8.055 3.415 ;
        RECT 1.055 1.98 7.95 2.24 ;
    END
  END virtpwr
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.55 7.945 2.67 ;
        RECT 5.72 1.55 6.37 2.67 ;
        RECT 4.165 1.55 4.815 2.67 ;
        RECT 2.61 1.55 3.26 2.67 ;
        RECT 1.055 1.55 1.705 2.67 ;
      LAYER met2 ;
        RECT 0.28 0 8.84 3.33 ;
      LAYER li ;
        RECT 1.055 1.55 7.95 1.81 ;
        RECT 1.055 2.41 7.95 2.67 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
END scs130lp_sleep_sergate_plv_21

MACRO scs130lp_sleep_sergate_plv_28
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sleep_sergate_plv_28 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 4.2 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.255 0.8 8.785 2.83 ;
    END
  END sleep
  PIN virtpwr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855 LAYER li ;
    ANTENNADIFFAREA 5.95 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
        RECT 6.51 1.105 7.155 3.575 ;
        RECT 4.955 1.105 5.58 3.575 ;
        RECT 3.4 1.105 4.025 3.575 ;
        RECT 1.845 1.105 2.47 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 1.055 2.84 8.055 3.415 ;
        RECT 1.055 1.12 7.95 1.38 ;
        RECT 1.055 1.98 7.95 2.24 ;
    END
  END virtpwr
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.55 7.945 2.67 ;
        RECT 5.72 1.55 6.37 2.67 ;
        RECT 4.165 1.55 4.815 2.67 ;
        RECT 2.61 1.55 3.26 2.67 ;
        RECT 1.055 1.55 1.705 2.67 ;
      LAYER met2 ;
        RECT 0.28 0 8.84 3.33 ;
      LAYER li ;
        RECT 1.055 1.55 7.95 1.81 ;
        RECT 1.055 2.41 7.95 2.67 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
END scs130lp_sleep_sergate_plv_28

MACRO scs130lp_srdlrtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_srdlrtp_1 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.105 1.08 0.435 1.41 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.045 1.09 5.635 1.42 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.555 1.815 11.915 3.075 ;
        RECT 11.745 0.255 11.915 3.075 ;
        RECT 11.555 0.255 11.915 1.135 ;
    END
  END Q
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.598 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.885 1.14 6.595 1.47 ;
    END
  END SLEEPB
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
      ANTENNAGATEAREA 0.472 LAYER met1 ;
      ANTENNAMAXAREACAR 1.399361 LAYER li ;
      ANTENNAMAXAREACAR 1.399361 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.886792 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.886792 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.181761 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 9.215 1.92 9.505 2.15 ;
        RECT 1.055 1.965 9.505 2.105 ;
        RECT 1.055 1.92 1.345 2.15 ;
      LAYER li ;
        RECT 9.225 1.55 9.955 2.15 ;
        RECT 0.945 1.92 1.315 2.255 ;
    END
  END RESETB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 11.93 2.945 ;
      LAYER li ;
        RECT 10.02 2.66 10.435 3.075 ;
        RECT 8.27 2.66 8.6 3.075 ;
        RECT 5.885 2.66 6.395 2.99 ;
        RECT 4.94 2.66 5.635 2.99 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12 0.085 ;
        RECT 11.125 -0.085 11.375 0.965 ;
        RECT 8.61 -0.085 8.94 0.365 ;
        RECT 6.15 -0.085 6.48 0.63 ;
        RECT 3.66 -0.085 3.99 0.355 ;
        RECT 0.945 -0.085 1.195 0.845 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
      LAYER li ;
        RECT 0 3.245 12 3.415 ;
        RECT 11.125 1.815 11.375 3.415 ;
        RECT 4.3 2.975 4.63 3.415 ;
        RECT 1.16 2.425 1.49 3.415 ;
        RECT 0.115 2.765 0.445 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 10.58 0.255 10.91 2.49 ;
      RECT 10.58 1.315 11.575 1.645 ;
      RECT 9.375 2.32 9.705 3.075 ;
      RECT 6.565 2.905 8.1 3.075 ;
      RECT 7.93 1.645 8.1 3.075 ;
      RECT 6.565 2.32 6.735 3.075 ;
      RECT 2.96 2.635 4.77 2.805 ;
      RECT 4.6 2.32 4.77 2.805 ;
      RECT 2.96 1.205 3.13 2.805 ;
      RECT 7.93 2.32 10.295 2.49 ;
      RECT 10.125 0.255 10.295 2.49 ;
      RECT 4.6 2.32 6.735 2.49 ;
      RECT 7.93 1.645 8.365 1.935 ;
      RECT 2.96 1.205 3.39 1.445 ;
      RECT 9.92 0.255 10.295 0.675 ;
      RECT 2.45 2.415 2.78 3.075 ;
      RECT 2.5 0.865 2.78 3.075 ;
      RECT 7.27 1.98 7.76 2.735 ;
      RECT 7.59 1.305 7.76 2.735 ;
      RECT 3.3 2.295 4.43 2.465 ;
      RECT 4.26 1.98 4.43 2.465 ;
      RECT 3.3 1.615 3.47 2.465 ;
      RECT 4.26 1.98 7.76 2.15 ;
      RECT 3.3 1.615 3.73 1.785 ;
      RECT 3.56 0.865 3.73 1.785 ;
      RECT 7.59 1.305 9.055 1.475 ;
      RECT 8.885 1.035 9.765 1.365 ;
      RECT 2.5 0.865 3.73 1.035 ;
      RECT 2.36 0.595 2.67 0.925 ;
      RECT 8.18 0.535 9.455 0.705 ;
      RECT 9.125 0.255 9.455 0.705 ;
      RECT 8.18 0.255 8.43 0.705 ;
      RECT 6.71 1.64 7.04 1.81 ;
      RECT 6.87 1.14 7.04 1.81 ;
      RECT 6.87 1.14 7.42 1.31 ;
      RECT 7.17 0.595 7.42 1.31 ;
      RECT 7.17 0.875 8.715 1.135 ;
      RECT 3.64 1.955 4.07 2.125 ;
      RECT 3.9 0.525 4.07 2.125 ;
      RECT 2 1.095 2.33 1.425 ;
      RECT 2 0.255 2.17 1.425 ;
      RECT 5.805 0.8 7 0.97 ;
      RECT 6.83 0.255 7 0.97 ;
      RECT 3.9 0.525 4.535 0.925 ;
      RECT 4.205 0.255 4.535 0.925 ;
      RECT 5.805 0.255 5.975 0.97 ;
      RECT 2.84 0.525 4.535 0.695 ;
      RECT 7.59 0.255 7.92 0.585 ;
      RECT 2.84 0.255 3.01 0.695 ;
      RECT 6.83 0.255 7.92 0.425 ;
      RECT 4.205 0.255 5.975 0.425 ;
      RECT 2 0.255 3.01 0.425 ;
      RECT 4.375 1.64 5.735 1.81 ;
      RECT 4.375 1.105 4.875 1.81 ;
      RECT 4.705 0.595 4.875 1.81 ;
      RECT 4.705 0.595 5.22 0.92 ;
      RECT 1.66 2.415 1.99 3.075 ;
      RECT 1.66 0.465 1.83 3.075 ;
      RECT 1.375 0.465 1.83 0.845 ;
      RECT 0.615 2.425 0.945 3.075 ;
      RECT 0.605 0.74 0.775 2.595 ;
      RECT 0.605 1.58 1.47 1.75 ;
      RECT 1.14 1.015 1.47 1.75 ;
      RECT 0.115 0.74 0.775 0.91 ;
      RECT 0.115 0.465 0.445 0.91 ;
  END
END scs130lp_srdlrtp_1

MACRO scs130lp_srdlstp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_srdlstp_1 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 0.955 0.455 1.78 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.285 1.48 8.615 2.15 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5943 LAYER li ;
    PORT
      LAYER li ;
        RECT 12.505 0.265 12.835 3.075 ;
    END
  END Q
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.409 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.435 0.255 5.765 0.56 ;
        RECT 5.435 0.255 5.635 0.67 ;
        RECT 1.98 0.255 5.765 0.425 ;
        RECT 1.98 0.255 2.31 0.475 ;
    END
  END SETB
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.598 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.685 1.48 11.055 2.15 ;
    END
  END SLEEPB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 12.89 2.945 ;
      LAYER li ;
        RECT 9.245 2.66 9.94 2.99 ;
        RECT 8.6 2.66 8.995 2.99 ;
        RECT 6.81 2.655 7.14 2.985 ;
        RECT 4.615 2.655 5.155 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 12.96 0.085 ;
        RECT 12.075 -0.085 12.325 1.145 ;
        RECT 11.055 -0.085 11.305 1.095 ;
        RECT 9.715 -0.085 10.045 1.31 ;
        RECT 6.82 -0.085 7.15 1.015 ;
        RECT 5.935 -0.085 6.185 0.945 ;
        RECT 1.835 0.645 2.165 1.31 ;
        RECT 1.64 0.645 2.165 0.815 ;
        RECT 1.64 -0.085 1.81 0.815 ;
        RECT 0.095 -0.085 0.345 0.785 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 12.96 3.415 ;
        RECT 12.005 1.815 12.335 3.415 ;
        RECT 1.61 2.845 1.94 3.415 ;
        RECT 0.64 2.32 0.97 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 11.31 1.475 11.64 2.495 ;
      RECT 11.485 1.315 12.335 1.645 ;
      RECT 11.485 0.635 11.815 1.645 ;
      RECT 8.05 2.745 8.43 3.075 ;
      RECT 8.26 2.32 8.43 3.075 ;
      RECT 10.255 0.635 10.505 2.86 ;
      RECT 8.26 2.32 10.505 2.49 ;
      RECT 10.255 0.635 10.595 1.095 ;
      RECT 3.185 2.905 4.4 3.075 ;
      RECT 4.23 1.125 4.4 3.075 ;
      RECT 3.185 1.765 3.355 3.075 ;
      RECT 4.23 2.315 8.09 2.485 ;
      RECT 7.92 1.14 8.09 2.485 ;
      RECT 9.065 1.14 9.395 2.15 ;
      RECT 3.025 1.765 3.355 2.095 ;
      RECT 4.07 1.125 4.4 1.455 ;
      RECT 7.92 1.14 9.395 1.31 ;
      RECT 8.425 0.85 8.755 1.31 ;
      RECT 4.64 1.975 7.75 2.145 ;
      RECT 7.58 0.8 7.75 2.145 ;
      RECT 7.42 1.685 7.75 2.145 ;
      RECT 4.64 1.625 4.97 2.145 ;
      RECT 7.58 0.8 8.205 0.97 ;
      RECT 7.875 0.34 8.205 0.97 ;
      RECT 3.59 2.075 3.92 2.735 ;
      RECT 3.67 0.595 3.84 2.735 ;
      RECT 5.56 1.455 5.89 1.805 ;
      RECT 5.14 1.455 7.25 1.625 ;
      RECT 7.08 1.185 7.41 1.515 ;
      RECT 4.57 1.285 5.31 1.455 ;
      RECT 4.57 0.595 4.74 1.455 ;
      RECT 3.67 0.595 4.74 0.895 ;
      RECT 5.48 1.115 6.64 1.285 ;
      RECT 6.39 0.615 6.64 1.285 ;
      RECT 5.48 0.84 5.65 1.285 ;
      RECT 5.015 0.84 5.65 1.01 ;
      RECT 5.015 0.595 5.265 1.01 ;
      RECT 2.685 2.265 3.015 3.075 ;
      RECT 1.15 1.98 1.4 2.86 ;
      RECT 1.15 2.505 3.015 2.675 ;
      RECT 1.3 0.63 1.47 2.675 ;
      RECT 2.685 1.425 2.855 3.075 ;
      RECT 2.685 1.425 3.5 1.595 ;
      RECT 3.33 0.595 3.5 1.595 ;
      RECT 1.045 0.63 1.47 1.31 ;
      RECT 2.88 0.595 3.5 0.815 ;
      RECT 2.145 1.48 2.515 2.335 ;
      RECT 2.345 0.85 2.515 2.335 ;
      RECT 2.345 0.985 3.16 1.255 ;
      RECT 2.345 0.85 2.69 1.255 ;
      RECT 0.105 1.98 0.435 2.66 ;
      RECT 0.105 1.98 0.855 2.15 ;
      RECT 0.685 0.325 0.855 2.15 ;
      RECT 0.685 1.48 1.13 1.81 ;
      RECT 0.525 0.325 0.855 0.785 ;
  END
END scs130lp_srdlstp_1

MACRO scs130lp_srdlxtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_srdlxtp_1 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.985 0.785 1.315 1.115 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.885 0.845 6.41 1.78 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 8.675 1.815 9.005 3.075 ;
        RECT 8.835 0.255 9.005 3.075 ;
        RECT 8.675 0.255 9.005 1.135 ;
    END
  END Q
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.015 0.775 7.555 1.41 ;
    END
  END SLEEPB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 9.05 2.945 ;
      LAYER li ;
        RECT 5.815 2.525 7.33 2.695 ;
        RECT 7 1.655 7.33 2.695 ;
        RECT 4.71 2.72 6.145 2.89 ;
        RECT 5.815 2.415 6.145 2.89 ;
        RECT 4.71 2.415 5.155 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.12 0.085 ;
        RECT 8.245 -0.085 8.495 1.135 ;
        RECT 7.14 -0.085 7.47 0.605 ;
        RECT 4.64 -0.085 4.97 0.675 ;
        RECT 1.825 -0.085 2.155 0.445 ;
        RECT 0.115 -0.085 0.365 1.335 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.12 3.415 ;
        RECT 8.175 1.815 8.505 3.415 ;
        RECT 1.61 2.775 1.94 3.415 ;
        RECT 0.115 2.395 0.365 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 7.63 1.815 7.96 2.495 ;
      RECT 7.79 0.255 7.96 2.495 ;
      RECT 7.79 1.315 8.665 1.645 ;
      RECT 7.79 0.255 8.03 1.645 ;
      RECT 7.7 0.255 8.03 0.605 ;
      RECT 2.31 2.905 4.375 3.075 ;
      RECT 4.205 1.185 4.375 3.075 ;
      RECT 3.15 1.965 3.475 3.075 ;
      RECT 2.31 1.625 2.48 3.075 ;
      RECT 6.58 0.505 6.83 2.335 ;
      RECT 4.205 2.075 6.83 2.245 ;
      RECT 2.31 1.625 2.64 1.955 ;
      RECT 0.875 1.625 1.205 1.955 ;
      RECT 0.875 1.625 2.64 1.795 ;
      RECT 4.045 1.185 4.375 1.515 ;
      RECT 5.99 0.505 6.83 0.675 ;
      RECT 5.99 0.255 6.32 0.675 ;
      RECT 4.585 1.575 5.615 1.905 ;
      RECT 5.445 0.255 5.615 1.905 ;
      RECT 5.43 0.255 5.76 0.675 ;
      RECT 3.69 2.075 4.02 2.735 ;
      RECT 3.69 0.845 3.86 2.735 ;
      RECT 4.945 0.845 5.275 1.175 ;
      RECT 3.46 0.845 5.275 1.015 ;
      RECT 3.46 0.255 3.79 1.015 ;
      RECT 2.65 2.445 2.98 2.735 ;
      RECT 2.81 1.625 2.98 2.735 ;
      RECT 2.81 1.625 3.29 1.795 ;
      RECT 3.12 0.505 3.29 1.795 ;
      RECT 2.36 0.505 3.29 0.675 ;
      RECT 2.36 0.255 2.69 0.675 ;
      RECT 0.535 2.395 0.875 3.075 ;
      RECT 0.535 0.875 0.705 3.075 ;
      RECT 0.535 1.285 2.95 1.455 ;
      RECT 2.62 1.055 2.95 1.455 ;
      RECT 0.535 0.875 0.795 1.455 ;
      RECT 1.86 0.615 2.19 1.095 ;
      RECT 1.485 0.615 2.19 0.785 ;
      RECT 1.165 0.255 1.655 0.615 ;
      RECT 1.11 2.435 1.44 3.075 ;
      RECT 1.11 2.435 2.105 2.605 ;
      RECT 1.775 1.965 2.105 2.605 ;
  END
END scs130lp_srdlxtp_1

MACRO scs130lp_sregrbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sregrbp_1 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.87 1.18 4.195 1.515 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.125 1.89 1.455 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.98 1.18 3.3 1.855 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.48 1.635 2.45 1.805 ;
        RECT 2.13 1.285 2.45 1.805 ;
        RECT 0.48 1.475 1.315 1.805 ;
    END
  END SCE
  PIN ASYNC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 1.071847 LAYER li ;
      ANTENNAMAXAREACAR 1.071847 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.995495 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.995495 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 11.135 1.92 11.425 2.15 ;
        RECT 7.775 1.965 11.425 2.105 ;
        RECT 7.775 1.92 8.065 2.15 ;
      LAYER li ;
        RECT 11.165 1.805 11.835 2.095 ;
        RECT 11.165 1.805 11.395 2.15 ;
        RECT 7.745 1.375 8.075 1.705 ;
        RECT 7.745 1.375 8.035 2.15 ;
    END
  END ASYNC
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    ANTENNADIFFAREA 0.5985 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 13.13 1.965 13.765 2.105 ;
        RECT 13.055 1.18 13.345 1.41 ;
        RECT 13.13 1.18 13.27 2.105 ;
      LAYER li ;
        RECT 12.965 0.265 13.325 2.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    ANTENNADIFFAREA 0.5985 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 14.015 1.92 14.305 2.15 ;
        RECT 14.09 1.225 14.23 2.15 ;
        RECT 13.595 1.225 14.23 1.365 ;
      LAYER li ;
        RECT 13.905 1.835 14.31 3.065 ;
        RECT 14.14 0.265 14.31 3.065 ;
        RECT 13.935 0.265 14.31 1.145 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 14.4 0.085 ;
        RECT 13.505 -0.085 13.755 1.145 ;
        RECT 12.005 -0.085 12.255 0.725 ;
        RECT 10.655 -0.085 10.985 0.805 ;
        RECT 8.635 -0.085 8.885 1.195 ;
        RECT 7.05 -0.085 7.38 1.195 ;
        RECT 4.335 -0.085 4.665 0.65 ;
        RECT 2.795 -0.085 3.045 0.675 ;
        RECT 1.105 -0.085 1.435 0.675 ;
        RECT 0.115 -0.085 0.365 0.71 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 14.4 3.415 ;
        RECT 13.395 2.675 13.725 3.415 ;
        RECT 11.71 2.275 12.04 3.415 ;
        RECT 10.69 2.68 11.02 3.415 ;
        RECT 8.7 1.885 9.03 3.415 ;
        RECT 7.595 2.68 7.925 3.415 ;
        RECT 6.57 2.295 6.82 3.415 ;
        RECT 4.215 2.045 4.545 3.415 ;
        RECT 2.645 2.845 2.975 3.415 ;
        RECT 0.865 2.635 1.195 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 9.215 1.55 9.505 1.78 ;
      RECT 5.375 1.55 5.665 1.78 ;
      RECT 5.375 1.595 9.505 1.735 ;
      RECT 5.375 0.44 5.665 0.67 ;
      RECT 3.455 0.44 3.745 0.67 ;
      RECT 3.455 0.485 5.665 0.625 ;
    LAYER li ;
      RECT 12.255 2.235 12.585 2.915 ;
      RECT 12.255 2.325 13.725 2.495 ;
      RECT 13.555 1.325 13.725 2.495 ;
      RECT 12.255 2.235 12.78 2.495 ;
      RECT 12.61 0.265 12.78 2.495 ;
      RECT 13.555 1.325 13.96 1.655 ;
      RECT 12.435 0.265 12.78 0.725 ;
      RECT 11.2 2.33 11.53 3.065 ;
      RECT 10.58 2.33 11.53 2.5 ;
      RECT 10.58 1.455 10.75 2.5 ;
      RECT 10.42 1.765 10.75 2.095 ;
      RECT 12.1 1.455 12.43 1.785 ;
      RECT 10.58 1.455 12.43 1.625 ;
      RECT 11.445 0.265 11.775 1.625 ;
      RECT 9.64 2.025 9.97 2.905 ;
      RECT 9.875 0.435 10.045 2.195 ;
      RECT 10.78 0.985 11.11 1.275 ;
      RECT 9.605 0.985 11.11 1.195 ;
      RECT 9.605 0.435 10.045 1.195 ;
      RECT 8.22 1.885 8.47 2.725 ;
      RECT 7.05 1.885 7.38 2.725 ;
      RECT 7.05 2.33 8.47 2.5 ;
      RECT 6.58 1.885 7.38 2.115 ;
      RECT 8.255 0.575 8.425 2.725 ;
      RECT 6.58 1.785 6.91 2.115 ;
      RECT 8.255 1.375 9.065 1.705 ;
      RECT 7.87 0.575 8.425 1.195 ;
      RECT 5.67 2.435 6.39 2.755 ;
      RECT 6.22 0.575 6.39 2.755 ;
      RECT 7.175 1.375 7.505 1.705 ;
      RECT 6.22 1.375 7.505 1.545 ;
      RECT 6.22 0.575 6.47 1.545 ;
      RECT 5.24 2.085 5.49 2.755 ;
      RECT 5.24 2.085 6.04 2.255 ;
      RECT 5.87 0.44 6.04 2.255 ;
      RECT 5.405 0.44 6.04 1.035 ;
      RECT 4.725 1.735 5.03 3.065 ;
      RECT 5.03 1.55 5.69 1.905 ;
      RECT 5.03 0.265 5.2 1.905 ;
      RECT 4.845 0.265 5.2 1.045 ;
      RECT 3.865 1.695 4.035 3.065 ;
      RECT 3.865 1.695 4.545 1.865 ;
      RECT 4.375 0.83 4.545 1.865 ;
      RECT 4.375 1.225 4.85 1.555 ;
      RECT 3.905 0.83 4.545 1 ;
      RECT 3.905 0.265 4.155 1 ;
      RECT 3.155 2.675 3.485 3.065 ;
      RECT 3.155 2.675 3.685 2.845 ;
      RECT 3.515 0.265 3.685 2.845 ;
      RECT 3.225 0.265 3.715 0.675 ;
      RECT 1.685 2.495 2.015 3.065 ;
      RECT 1.685 2.495 2.8 2.665 ;
      RECT 2.63 0.855 2.8 2.665 ;
      RECT 2.63 2.165 3.335 2.495 ;
      RECT 2.135 0.855 2.8 1.025 ;
      RECT 2.135 0.265 2.305 1.025 ;
      RECT 1.975 0.265 2.305 0.675 ;
      RECT 0.13 2.635 0.685 3.065 ;
      RECT 0.13 0.89 0.3 3.065 ;
      RECT 0.13 1.985 2.28 2.315 ;
      RECT 0.13 0.89 1.14 1.22 ;
      RECT 0.545 0.265 0.875 1.22 ;
      RECT 9.245 1.375 9.695 1.78 ;
  END
END scs130lp_sregrbp_1

MACRO scs130lp_sregsbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_sregsbp_1 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.87 1.18 4.195 1.515 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.56 1.125 1.89 1.455 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.126 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.98 1.18 3.3 1.855 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.48 1.635 2.45 1.805 ;
        RECT 2.13 1.285 2.45 1.805 ;
        RECT 0.48 1.475 1.315 1.805 ;
    END
  END SCE
  PIN ASYNC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
      ANTENNAGATEAREA 0.444 LAYER met1 ;
      ANTENNAMAXAREACAR 1.071847 LAYER li ;
      ANTENNAMAXAREACAR 1.071847 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.995495 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.995495 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.13018 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 11.135 1.92 11.425 2.15 ;
        RECT 7.775 1.965 11.425 2.105 ;
        RECT 7.775 1.92 8.065 2.15 ;
      LAYER li ;
        RECT 11.165 1.805 11.835 2.095 ;
        RECT 11.165 1.805 11.395 2.15 ;
        RECT 7.745 1.375 8.075 1.705 ;
        RECT 7.745 1.375 8.035 2.15 ;
    END
  END ASYNC
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    ANTENNADIFFAREA 0.5985 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 14.015 1.92 14.305 2.15 ;
        RECT 14.09 1.295 14.23 2.15 ;
        RECT 13.595 1.965 14.305 2.105 ;
      LAYER li ;
        RECT 13.905 1.835 14.31 3.065 ;
        RECT 14.14 0.265 14.31 3.065 ;
        RECT 13.935 0.265 14.31 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    ANTENNADIFFAREA 0.5985 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 13.055 1.225 13.765 1.365 ;
        RECT 13.055 1.18 13.345 1.41 ;
        RECT 13.13 1.18 13.27 2.035 ;
      LAYER li ;
        RECT 12.965 0.265 13.325 2.145 ;
    END
  END QN
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
      LAYER li ;
        RECT 0 -0.085 14.4 0.085 ;
        RECT 13.505 -0.085 13.755 1.145 ;
        RECT 12.005 -0.085 12.255 0.725 ;
        RECT 10.655 -0.085 10.985 0.805 ;
        RECT 8.635 -0.085 8.885 1.195 ;
        RECT 7.05 -0.085 7.38 1.195 ;
        RECT 4.335 -0.085 4.665 0.65 ;
        RECT 2.795 -0.085 3.045 0.675 ;
        RECT 1.105 -0.085 1.435 0.675 ;
        RECT 0.115 -0.085 0.365 0.71 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
      LAYER li ;
        RECT 0 3.245 14.4 3.415 ;
        RECT 13.395 2.675 13.725 3.415 ;
        RECT 11.71 2.275 12.04 3.415 ;
        RECT 10.69 2.68 11.02 3.415 ;
        RECT 8.7 1.885 9.03 3.415 ;
        RECT 7.595 2.68 7.925 3.415 ;
        RECT 6.57 2.295 6.82 3.415 ;
        RECT 4.215 2.045 4.545 3.415 ;
        RECT 2.645 2.845 2.975 3.415 ;
        RECT 0.865 2.635 1.195 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 9.215 1.55 9.505 1.78 ;
      RECT 5.375 1.55 5.665 1.78 ;
      RECT 5.375 1.595 9.505 1.735 ;
      RECT 5.375 0.44 5.665 0.67 ;
      RECT 2.015 0.44 2.305 0.67 ;
      RECT 2.015 0.485 5.665 0.625 ;
    LAYER li ;
      RECT 12.255 2.235 12.585 2.915 ;
      RECT 12.255 2.325 13.725 2.495 ;
      RECT 13.555 1.325 13.725 2.495 ;
      RECT 12.255 2.235 12.78 2.495 ;
      RECT 12.61 0.265 12.78 2.495 ;
      RECT 13.555 1.325 13.96 1.655 ;
      RECT 12.435 0.265 12.78 0.725 ;
      RECT 11.2 2.33 11.53 3.065 ;
      RECT 10.58 2.33 11.53 2.5 ;
      RECT 10.58 1.455 10.75 2.5 ;
      RECT 10.42 1.765 10.75 2.095 ;
      RECT 12.1 1.455 12.43 1.785 ;
      RECT 10.58 1.455 12.43 1.625 ;
      RECT 11.445 0.265 11.775 1.625 ;
      RECT 9.64 2.025 9.97 2.905 ;
      RECT 9.875 0.435 10.045 2.195 ;
      RECT 10.78 0.985 11.11 1.275 ;
      RECT 9.605 0.985 11.11 1.195 ;
      RECT 9.605 0.435 10.045 1.195 ;
      RECT 8.22 1.885 8.47 2.725 ;
      RECT 7.05 1.885 7.38 2.725 ;
      RECT 7.05 2.33 8.47 2.5 ;
      RECT 6.58 1.885 7.38 2.115 ;
      RECT 8.255 0.575 8.425 2.725 ;
      RECT 6.58 1.785 6.91 2.115 ;
      RECT 8.255 1.375 9.065 1.705 ;
      RECT 7.87 0.575 8.425 1.195 ;
      RECT 5.67 2.435 6.39 2.755 ;
      RECT 6.22 0.575 6.39 2.755 ;
      RECT 7.175 1.375 7.505 1.705 ;
      RECT 6.22 1.375 7.505 1.545 ;
      RECT 6.22 0.575 6.47 1.545 ;
      RECT 5.24 2.085 5.49 2.755 ;
      RECT 5.24 2.085 6.04 2.255 ;
      RECT 5.87 0.44 6.04 2.255 ;
      RECT 5.405 0.44 6.04 1.035 ;
      RECT 4.725 1.735 5.03 3.065 ;
      RECT 5.03 1.55 5.69 1.905 ;
      RECT 5.03 0.265 5.2 1.905 ;
      RECT 4.845 0.265 5.2 1.045 ;
      RECT 3.865 1.695 4.035 3.065 ;
      RECT 3.865 1.695 4.545 1.865 ;
      RECT 4.375 0.83 4.545 1.865 ;
      RECT 4.375 1.225 4.85 1.555 ;
      RECT 3.905 0.83 4.545 1 ;
      RECT 3.905 0.265 4.155 1 ;
      RECT 3.155 2.675 3.485 3.065 ;
      RECT 3.155 2.675 3.685 2.845 ;
      RECT 3.515 0.265 3.685 2.845 ;
      RECT 3.225 0.265 3.715 0.675 ;
      RECT 1.685 2.495 2.015 3.065 ;
      RECT 1.685 2.495 2.8 2.665 ;
      RECT 2.63 0.855 2.8 2.665 ;
      RECT 2.63 2.165 3.335 2.495 ;
      RECT 2.135 0.855 2.8 1.025 ;
      RECT 2.135 0.265 2.305 1.025 ;
      RECT 1.975 0.265 2.305 0.675 ;
      RECT 0.13 2.635 0.685 3.065 ;
      RECT 0.13 0.89 0.3 3.065 ;
      RECT 0.13 1.985 2.28 2.315 ;
      RECT 0.13 0.89 1.14 1.22 ;
      RECT 0.545 0.265 0.875 1.22 ;
      RECT 9.245 1.375 9.695 1.78 ;
  END
END scs130lp_sregsbp_1

MACRO scs130lp_srsdfrtn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_srsdfrtn_1 0 0 ;
  SIZE 18.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.205 1.555 10.685 1.84 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.18 1.805 1.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5859 LAYER li ;
    PORT
      LAYER li ;
        RECT 17.795 0.265 18.135 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.598 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.9 1.61 8.14 1.78 ;
        RECT 7.805 1.215 8.14 1.78 ;
        RECT 6.9 0.255 7.07 1.78 ;
        RECT 4.605 0.255 7.07 0.425 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.605 2.87 2.275 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.585 1.095 0.915 1.78 ;
    END
  END SCE
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.598 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.195 1.295 11.56 1.78 ;
    END
  END SLEEPB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 18.17 2.945 ;
        RECT 11.615 2.66 11.905 2.945 ;
        RECT 8.255 2.66 8.545 2.945 ;
        RECT 7.775 2.66 8.065 2.945 ;
      LAYER li ;
        RECT 10.845 2.905 12.05 3.075 ;
        RECT 11.645 2.29 12.05 3.075 ;
        RECT 10.845 2.35 11.015 3.075 ;
        RECT 8.285 2.69 9.24 3.02 ;
        RECT 7.415 2.69 8.035 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 18.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 18.24 0.085 ;
        RECT 17.365 -0.085 17.615 1.145 ;
        RECT 15.12 -0.085 15.45 0.935 ;
        RECT 11.91 -0.085 12.16 0.445 ;
        RECT 8.825 -0.085 9.075 0.675 ;
        RECT 7.78 -0.085 8.11 0.365 ;
        RECT 3.835 -0.085 4.165 0.755 ;
        RECT 0.535 -0.085 0.865 0.715 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 18.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 18.24 3.415 ;
        RECT 17.375 1.815 17.625 3.415 ;
        RECT 16.385 2.295 16.635 3.415 ;
        RECT 15.445 2.305 15.695 3.415 ;
        RECT 4.285 2.075 4.455 3.415 ;
        RECT 2.67 2.785 2.92 3.415 ;
        RECT 0.78 2.435 1.11 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 14.015 1.92 14.305 2.15 ;
      RECT 6.335 1.92 6.625 2.15 ;
      RECT 3.455 1.92 3.745 2.15 ;
      RECT 3.455 1.965 14.305 2.105 ;
    LAYER li ;
      RECT 16.84 2.435 17.17 3.075 ;
      RECT 16.98 1.315 17.17 3.075 ;
      RECT 16.98 1.315 17.625 1.645 ;
      RECT 16.98 0.265 17.15 3.075 ;
      RECT 16.82 0.265 17.15 0.725 ;
      RECT 13.655 2.565 14.925 2.735 ;
      RECT 14.755 1.965 14.925 2.735 ;
      RECT 13.655 0.785 13.905 2.735 ;
      RECT 14.87 1.105 15.04 2.135 ;
      RECT 16.48 0.895 16.81 1.565 ;
      RECT 14.87 1.105 15.79 1.275 ;
      RECT 15.62 0.255 15.79 1.275 ;
      RECT 13.825 0.595 14.155 0.955 ;
      RECT 16.48 0.255 16.65 1.565 ;
      RECT 15.62 0.255 16.65 0.425 ;
      RECT 15.875 1.805 16.205 2.755 ;
      RECT 16.035 0.595 16.205 2.755 ;
      RECT 15.21 1.805 16.205 2.135 ;
      RECT 16.035 0.595 16.305 0.935 ;
      RECT 12.77 2.905 15.265 3.075 ;
      RECT 15.095 2.305 15.265 3.075 ;
      RECT 12.77 2.245 13.1 3.075 ;
      RECT 14.415 1.625 14.585 2.395 ;
      RECT 8.355 1.67 9.96 1.84 ;
      RECT 9.63 1.59 9.96 1.84 ;
      RECT 14.53 0.255 14.7 1.795 ;
      RECT 8.355 0.875 8.525 1.84 ;
      RECT 7.24 0.875 7.57 1.44 ;
      RECT 7.24 0.875 9.865 1.045 ;
      RECT 9.535 0.255 9.865 1.045 ;
      RECT 11.535 0.615 12.595 0.785 ;
      RECT 12.425 0.255 12.595 0.785 ;
      RECT 13.325 0.255 13.655 0.615 ;
      RECT 11.535 0.255 11.705 0.785 ;
      RECT 12.425 0.255 14.7 0.425 ;
      RECT 9.535 0.255 11.705 0.425 ;
      RECT 14.075 1.125 14.245 2.15 ;
      RECT 14.075 1.125 14.36 1.455 ;
      RECT 12.25 1.715 12.58 2.755 ;
      RECT 12.25 1.905 13.485 2.075 ;
      RECT 13.315 0.955 13.485 2.075 ;
      RECT 8.695 1.215 9.025 1.5 ;
      RECT 8.695 1.215 10.205 1.385 ;
      RECT 10.035 0.595 10.205 1.385 ;
      RECT 11.195 0.955 13.485 1.125 ;
      RECT 12.765 0.595 13.095 1.125 ;
      RECT 11.195 0.595 11.365 1.125 ;
      RECT 10.035 0.595 11.365 0.765 ;
      RECT 5.21 2.905 7.245 3.075 ;
      RECT 7.075 2.35 7.245 3.075 ;
      RECT 5.21 1.605 5.38 3.075 ;
      RECT 9.41 2.725 10.675 2.895 ;
      RECT 10.505 2.01 10.675 2.895 ;
      RECT 11.195 1.95 11.445 2.735 ;
      RECT 9.41 2.35 9.58 2.895 ;
      RECT 7.075 2.35 9.58 2.52 ;
      RECT 10.505 2.01 11.445 2.18 ;
      RECT 11.91 1.375 12.08 2.12 ;
      RECT 11.195 1.95 12.08 2.12 ;
      RECT 10.855 0.935 11.025 2.18 ;
      RECT 5.05 1.605 5.38 1.935 ;
      RECT 12.75 1.375 13.145 1.735 ;
      RECT 11.91 1.375 13.145 1.545 ;
      RECT 10.42 0.935 11.025 1.265 ;
      RECT 5.55 1.275 5.985 2.735 ;
      RECT 10.08 2.01 10.335 2.555 ;
      RECT 5.55 2.32 6.905 2.49 ;
      RECT 6.735 1.95 6.905 2.49 ;
      RECT 6.735 2.01 10.335 2.18 ;
      RECT 6.735 1.95 8.185 2.18 ;
      RECT 7.24 0.535 8.645 0.705 ;
      RECT 8.315 0.255 8.645 0.705 ;
      RECT 7.24 0.365 7.57 0.705 ;
      RECT 3.09 2.905 4.115 3.075 ;
      RECT 3.945 1.735 4.115 3.075 ;
      RECT 1.6 2.445 1.93 3.075 ;
      RECT 3.09 2.445 3.26 3.075 ;
      RECT 4.635 2.105 4.965 2.755 ;
      RECT 1.6 2.445 3.26 2.615 ;
      RECT 3.04 1.265 3.21 2.615 ;
      RECT 4.635 1.265 4.805 2.755 ;
      RECT 3.945 1.735 4.805 1.905 ;
      RECT 6.34 0.935 6.67 1.435 ;
      RECT 4.635 1.265 5.38 1.435 ;
      RECT 5.21 0.935 5.38 1.435 ;
      RECT 1.975 1.265 3.21 1.435 ;
      RECT 1.975 0.595 2.145 1.435 ;
      RECT 5.21 0.935 6.67 1.105 ;
      RECT 1.5 0.595 2.145 0.925 ;
      RECT 2.4 0.925 4.7 1.095 ;
      RECT 4.37 0.595 4.7 1.095 ;
      RECT 2.4 0.595 2.57 1.095 ;
      RECT 3.485 1.265 3.735 2.735 ;
      RECT 3.38 1.265 3.735 1.595 ;
      RECT 1.07 0.255 1.32 0.925 ;
      RECT 2.75 0.255 3.08 0.755 ;
      RECT 1.07 0.255 3.08 0.425 ;
      RECT 0.105 1.95 0.61 3.075 ;
      RECT 1.975 1.945 2.305 2.275 ;
      RECT 0.105 1.95 2.305 2.12 ;
      RECT 0.105 0.255 0.355 3.075 ;
      RECT 5.015 0.595 6.73 0.765 ;
      RECT 6.155 1.605 6.565 2.15 ;
  END
END scs130lp_srsdfrtn_1

MACRO scs130lp_srsdfrtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_srsdfrtp_1 0 0 ;
  SIZE 20.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 16.59 1.46 17.155 1.79 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.565 1.84 2.135 2.17 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5901 LAYER li ;
    PORT
      LAYER li ;
        RECT 20.205 0.265 20.535 2.15 ;
        RECT 19.995 1.815 20.325 3.075 ;
    END
  END Q
  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.598 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.92 1.55 4.25 1.88 ;
    END
  END RESETB
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.35 1.55 3.715 1.88 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.605 1.5 0.935 2.17 ;
    END
  END SCE
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.598 LAYER li ;
    PORT
      LAYER li ;
        RECT 18.235 1.12 18.565 1.45 ;
    END
  END SLEEPB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 20.57 2.945 ;
      LAYER li ;
        RECT 16.925 2.69 17.73 3.025 ;
        RECT 16.28 2.69 16.675 2.97 ;
        RECT 14.525 2.69 14.975 2.97 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 20.64 0.245 ;
      LAYER li ;
        RECT 0 -0.085 20.64 0.085 ;
        RECT 19.855 -0.085 20.025 1.145 ;
        RECT 18.805 -0.085 19.055 0.805 ;
        RECT 17.475 -0.085 17.805 0.61 ;
        RECT 13.125 -0.085 13.455 0.81 ;
        RECT 11.365 -0.085 11.695 0.985 ;
        RECT 8.02 -0.085 8.35 0.825 ;
        RECT 7.05 -0.085 7.38 0.835 ;
        RECT 3.615 -0.085 3.865 1.04 ;
        RECT 0.535 -0.085 0.865 0.99 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 20.64 3.575 ;
      LAYER li ;
        RECT 0 3.245 20.64 3.415 ;
        RECT 19.495 1.815 19.825 3.415 ;
        RECT 7.85 2.605 8.18 3.415 ;
        RECT 6.12 2.77 6.45 3.415 ;
        RECT 3.245 2.44 3.575 3.415 ;
        RECT 0.62 2.34 0.95 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 18.735 1.815 18.985 2.18 ;
      RECT 18.735 0.975 18.905 2.18 ;
      RECT 19.515 1.315 20.02 1.645 ;
      RECT 19.515 0.345 19.685 1.645 ;
      RECT 18.735 0.975 19.685 1.145 ;
      RECT 19.235 0.345 19.685 1.145 ;
      RECT 13.625 2.35 13.955 2.97 ;
      RECT 9.89 2.565 12.54 2.735 ;
      RECT 12.21 2.35 12.54 2.735 ;
      RECT 9.89 2.04 10.5 2.735 ;
      RECT 10.19 0.605 10.5 2.735 ;
      RECT 12.21 2.35 19.325 2.52 ;
      RECT 19.155 1.315 19.325 2.52 ;
      RECT 16.25 1.41 16.42 2.52 ;
      RECT 15.985 1.41 16.42 1.74 ;
      RECT 19.075 1.315 19.345 1.645 ;
      RECT 17.895 1.85 18.49 2.18 ;
      RECT 17.895 0.78 18.065 2.18 ;
      RECT 12.93 1.32 14.185 1.5 ;
      RECT 14.015 0.6 14.185 1.5 ;
      RECT 16.93 0.78 18.345 0.95 ;
      RECT 18.015 0.345 18.345 0.95 ;
      RECT 16.93 0.255 17.1 0.95 ;
      RECT 14.015 0.6 15.315 0.77 ;
      RECT 14.985 0.255 15.315 0.77 ;
      RECT 14.985 0.255 17.1 0.425 ;
      RECT 16.855 2.01 17.495 2.18 ;
      RECT 17.325 1.12 17.495 2.18 ;
      RECT 11.64 1.67 14.525 1.84 ;
      RECT 14.355 0.94 14.525 1.84 ;
      RECT 11.64 1.51 11.97 1.84 ;
      RECT 16.59 1.12 17.495 1.29 ;
      RECT 16.105 0.95 16.76 1.12 ;
      RECT 14.355 0.94 16.435 1.11 ;
      RECT 16.105 0.595 16.435 1.12 ;
      RECT 15.645 1.93 16.08 2.18 ;
      RECT 11.1 2.01 14.955 2.18 ;
      RECT 14.695 1.28 14.955 2.18 ;
      RECT 11.1 1.155 11.43 2.18 ;
      RECT 15.645 1.44 15.815 2.18 ;
      RECT 14.695 1.44 15.815 1.61 ;
      RECT 11.1 1.155 12.235 1.325 ;
      RECT 11.905 0.575 12.235 1.325 ;
      RECT 12.695 0.98 13.845 1.15 ;
      RECT 13.675 0.575 13.845 1.15 ;
      RECT 12.695 0.575 12.945 1.15 ;
      RECT 8.555 2.905 13.455 3.075 ;
      RECT 13.125 2.745 13.455 3.075 ;
      RECT 8.555 1.335 8.725 3.075 ;
      RECT 8.395 1.335 8.725 2.825 ;
      RECT 4.925 2.6 5.95 2.77 ;
      RECT 5.78 2.43 7.68 2.6 ;
      RECT 4.925 1.59 5.095 2.77 ;
      RECT 7.51 2.265 8.725 2.435 ;
      RECT 4.885 1.59 5.215 1.92 ;
      RECT 9.21 1.495 9.54 1.825 ;
      RECT 8.395 1.495 9.54 1.665 ;
      RECT 8.395 1.335 8.99 1.665 ;
      RECT 10.68 0.265 10.93 2.395 ;
      RECT 7.34 1.845 8.135 2.095 ;
      RECT 7.965 0.995 8.135 2.095 ;
      RECT 5.96 1.435 6.29 1.825 ;
      RECT 6.28 1.005 6.61 1.605 ;
      RECT 9.2 0.265 9.53 1.285 ;
      RECT 6.28 1.005 8.135 1.175 ;
      RECT 7.59 0.995 9.53 1.165 ;
      RECT 7.59 0.575 7.84 1.175 ;
      RECT 9.2 0.265 10.93 0.435 ;
      RECT 5.265 2.09 5.555 2.43 ;
      RECT 5.385 0.935 5.555 2.43 ;
      RECT 5.265 2.09 7.11 2.26 ;
      RECT 6.78 1.345 7.11 2.26 ;
      RECT 6.78 1.345 7.795 1.675 ;
      RECT 5.375 0.935 5.555 1.265 ;
      RECT 4.615 0.255 4.865 1.08 ;
      RECT 6.26 0.255 6.59 0.835 ;
      RECT 4.615 0.255 6.59 0.425 ;
      RECT 4.425 2.1 4.755 2.99 ;
      RECT 2.305 2.1 2.635 2.99 ;
      RECT 1.225 2.34 2.635 2.51 ;
      RECT 1.225 1.5 1.395 2.51 ;
      RECT 2.305 2.1 4.755 2.27 ;
      RECT 4.545 1.25 4.715 2.99 ;
      RECT 1.225 1.5 2.08 1.67 ;
      RECT 1.83 0.935 2.08 1.67 ;
      RECT 4.545 1.25 5.205 1.42 ;
      RECT 5.035 0.595 5.205 1.42 ;
      RECT 5.725 0.595 6.055 1.265 ;
      RECT 5.035 0.595 6.055 0.765 ;
      RECT 2.645 1.21 4.375 1.38 ;
      RECT 4.045 0.58 4.375 1.38 ;
      RECT 2.645 0.74 2.975 1.38 ;
      RECT 3.155 0.255 3.405 1.04 ;
      RECT 1.07 0.255 1.32 0.99 ;
      RECT 1.07 0.255 3.405 0.425 ;
      RECT 0.105 1.16 0.435 2.99 ;
      RECT 2.305 1.6 2.88 1.93 ;
      RECT 2.305 0.595 2.475 1.93 ;
      RECT 0.105 1.16 1.66 1.33 ;
      RECT 1.49 0.595 1.66 1.33 ;
      RECT 0.105 0.53 0.355 2.99 ;
      RECT 1.49 0.595 2.475 0.765 ;
  END
END scs130lp_srsdfrtp_1

MACRO scs130lp_srsdfstp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_srsdfstp_1 0 0 ;
  SIZE 18.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 14.965 1.18 15.235 2.15 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.545 1.43 1.875 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5733 LAYER li ;
    PORT
      LAYER li ;
        RECT 18.365 0.255 18.62 3.075 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.125 1.205 0.835 1.875 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.725 1.18 3.235 1.555 ;
    END
  END SCE
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.439 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.5 1.58 13.83 1.84 ;
    END
  END SETB
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.598 LAYER li ;
    PORT
      LAYER li ;
        RECT 15.935 1.22 16.26 2.15 ;
    END
  END SLEEPB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 18.65 2.945 ;
      LAYER li ;
        RECT 15.965 2.66 16.305 2.94 ;
        RECT 12.655 2.905 15.235 3.075 ;
        RECT 14.905 2.66 15.235 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 18.72 0.245 ;
      LAYER li ;
        RECT 0 -0.085 18.72 0.085 ;
        RECT 17.86 -0.085 18.19 1.015 ;
        RECT 16.085 -0.085 16.335 0.71 ;
        RECT 11.745 -0.085 11.995 0.955 ;
        RECT 10.775 -0.085 11.025 1.035 ;
        RECT 7.115 -0.085 7.365 0.96 ;
        RECT 5.465 -0.085 5.795 0.505 ;
        RECT 2.92 -0.085 3.25 1.01 ;
        RECT 1.94 -0.085 2.19 1.035 ;
        RECT 0.1 -0.085 0.43 1.035 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 18.72 3.575 ;
      LAYER li ;
        RECT 0 3.245 18.72 3.415 ;
        RECT 17.855 1.815 18.185 3.415 ;
        RECT 7.25 2.265 7.58 3.415 ;
        RECT 6.025 2.655 6.355 3.415 ;
        RECT 2.92 2.565 3.25 3.415 ;
        RECT 0.6 2.385 0.85 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 17.39 1.995 17.675 2.675 ;
      RECT 17.505 0.295 17.675 2.675 ;
      RECT 17.505 1.185 18.195 1.515 ;
      RECT 17.325 0.295 17.675 0.675 ;
      RECT 8.94 2.745 12.485 3.075 ;
      RECT 12.315 2.565 12.485 3.075 ;
      RECT 8.925 0.935 9.095 2.745 ;
      RECT 8.895 2.235 9.145 2.745 ;
      RECT 12.315 2.565 14.13 2.735 ;
      RECT 13.8 2.35 14.13 2.735 ;
      RECT 13.8 2.35 14.595 2.52 ;
      RECT 17.05 1.495 17.22 2.49 ;
      RECT 14.425 2.32 17.22 2.49 ;
      RECT 17.005 1.495 17.335 1.825 ;
      RECT 8.865 0.935 9.195 1.225 ;
      RECT 16.455 0.88 16.835 2.15 ;
      RECT 11.625 1.125 12.335 1.375 ;
      RECT 12.165 0.255 12.335 1.375 ;
      RECT 15.745 0.88 16.835 1.05 ;
      RECT 16.665 0.63 16.835 2.15 ;
      RECT 15.745 0.255 15.915 1.05 ;
      RECT 16.795 0.42 17.125 0.8 ;
      RECT 13.525 0.255 13.855 0.73 ;
      RECT 12.165 0.255 15.915 0.425 ;
      RECT 15.405 1.9 15.765 2.15 ;
      RECT 10.165 1.545 10.415 2.145 ;
      RECT 15.405 0.595 15.575 2.15 ;
      RECT 10.085 1.545 12.675 1.715 ;
      RECT 12.505 0.595 12.675 1.715 ;
      RECT 10.085 0.255 10.255 1.715 ;
      RECT 5.45 0.675 5.78 1.375 ;
      RECT 6.725 1.13 7.705 1.3 ;
      RECT 7.535 0.255 7.705 1.3 ;
      RECT 6.725 0.255 6.895 1.3 ;
      RECT 13.185 0.9 14.255 1.07 ;
      RECT 14.085 0.595 14.255 1.07 ;
      RECT 13.185 0.595 13.355 1.07 ;
      RECT 14.085 0.595 15.575 0.845 ;
      RECT 5.45 0.675 6.135 0.845 ;
      RECT 5.965 0.255 6.135 0.845 ;
      RECT 12.505 0.595 13.355 0.765 ;
      RECT 7.535 0.255 10.255 0.425 ;
      RECT 5.965 0.255 6.895 0.425 ;
      RECT 11.475 1.885 11.805 2.235 ;
      RECT 10.655 1.885 10.985 2.215 ;
      RECT 10.655 1.885 13.015 2.055 ;
      RECT 12.845 0.935 13.015 2.055 ;
      RECT 12.845 1.24 14.755 1.41 ;
      RECT 14.425 1.04 14.755 1.41 ;
      RECT 7.755 2.905 8.695 3.075 ;
      RECT 8.525 0.595 8.695 3.075 ;
      RECT 7.845 1.47 8.015 3.075 ;
      RECT 9.315 2.405 12.145 2.575 ;
      RECT 11.975 2.225 12.145 2.575 ;
      RECT 9.315 1.885 9.485 2.575 ;
      RECT 11.975 2.225 13.355 2.395 ;
      RECT 13.185 2.01 13.355 2.395 ;
      RECT 4.005 1.725 4.26 2.395 ;
      RECT 13.185 2.01 14.21 2.18 ;
      RECT 14.04 1.58 14.21 2.18 ;
      RECT 9.365 0.595 9.535 2.135 ;
      RECT 3.42 1.725 4.26 2.055 ;
      RECT 14.04 1.58 14.37 1.91 ;
      RECT 8.525 1.41 8.755 1.74 ;
      RECT 3.42 0.255 3.75 2.055 ;
      RECT 5.11 1.545 6.12 1.715 ;
      RECT 5.95 1.47 8.015 1.64 ;
      RECT 5.11 0.255 5.28 1.715 ;
      RECT 8.525 0.595 9.535 0.765 ;
      RECT 3.42 0.255 4.015 0.585 ;
      RECT 3.42 0.255 5.28 0.425 ;
      RECT 10.425 1.205 11.455 1.375 ;
      RECT 11.205 0.605 11.455 1.375 ;
      RECT 10.425 0.605 10.595 1.375 ;
      RECT 8.185 1.095 8.355 2.565 ;
      RECT 7.875 1.095 8.355 1.265 ;
      RECT 7.875 0.595 8.145 1.265 ;
      RECT 5.205 1.905 5.535 3.075 ;
      RECT 6.44 1.81 7.675 2.095 ;
      RECT 4.77 1.905 7.675 2.075 ;
      RECT 4.77 0.675 4.94 2.075 ;
      RECT 4.41 0.675 4.94 1.135 ;
      RECT 6.68 2.265 7.01 2.695 ;
      RECT 5.9 2.265 7.01 2.485 ;
      RECT 5.9 2.245 6.23 2.485 ;
      RECT 5.99 1.015 6.555 1.3 ;
      RECT 6.305 0.595 6.555 1.3 ;
      RECT 4.6 2.655 5.035 3.075 ;
      RECT 3.665 2.655 5.035 2.825 ;
      RECT 4.43 1.385 4.6 2.825 ;
      RECT 1.43 2.225 1.77 2.735 ;
      RECT 1.6 0.865 1.77 2.735 ;
      RECT 3.665 2.225 3.835 2.825 ;
      RECT 1.43 2.225 3.835 2.395 ;
      RECT 3.98 1.385 4.6 1.555 ;
      RECT 3.98 0.755 4.23 1.555 ;
      RECT 0.92 0.865 1.77 1.035 ;
      RECT 0.92 0.575 1.25 1.035 ;
      RECT 1.94 1.725 2.72 2.055 ;
      RECT 1.94 1.305 2.555 2.055 ;
      RECT 2.385 0.675 2.555 2.055 ;
      RECT 2.385 0.675 2.74 1.01 ;
      RECT 1.02 2.905 2.19 3.075 ;
      RECT 1.94 2.565 2.19 3.075 ;
      RECT 0.1 2.045 0.43 3.065 ;
      RECT 1.02 2.045 1.19 3.075 ;
      RECT 0.1 2.045 1.19 2.215 ;
  END
END scs130lp_srsdfstp_1

MACRO scs130lp_srsdfxtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_srsdfxtp_1 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.725 1.5 11.01 1.83 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.18 1.59 1.51 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 13.475 1.815 13.835 3.075 ;
        RECT 13.665 0.265 13.835 3.075 ;
        RECT 13.475 0.265 13.835 1.145 ;
    END
  END Q
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.159 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.075 1.75 2.49 2.15 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.795 1.18 2.275 1.51 ;
        RECT 1.795 0.84 1.965 1.51 ;
        RECT 0.585 0.84 1.965 1.01 ;
        RECT 0.425 0.985 0.755 1.315 ;
    END
  END SCE
  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.222 LAYER li ;
    PORT
      LAYER li ;
        RECT 11.52 0.255 11.85 0.65 ;
        RECT 9.805 0.255 11.85 0.425 ;
        RECT 9.805 0.255 10.135 0.575 ;
    END
  END SLEEPB
  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 13.85 2.945 ;
      LAYER li ;
        RECT 11.195 2.68 11.365 3.075 ;
        RECT 9.725 2.68 10.005 3.075 ;
    END
  END kapwr
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
      LAYER li ;
        RECT 0 -0.085 13.92 0.085 ;
        RECT 13.045 -0.085 13.295 1.145 ;
        RECT 12.02 -0.085 12.27 1.33 ;
        RECT 7.95 -0.085 8.28 0.915 ;
        RECT 4.805 -0.085 5.055 0.445 ;
        RECT 2.475 -0.085 2.645 0.67 ;
        RECT 0.595 -0.085 0.925 0.67 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
      LAYER li ;
        RECT 0 3.245 13.92 3.415 ;
        RECT 13.045 1.815 13.295 3.415 ;
        RECT 5.495 2.965 5.825 3.415 ;
        RECT 2.4 2.66 2.65 3.415 ;
        RECT 0.565 2.365 0.895 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 12.5 0.265 12.83 2.495 ;
      RECT 12.5 1.315 13.495 1.645 ;
      RECT 11.535 2.745 12.595 3.075 ;
      RECT 10.175 2.905 11.025 3.075 ;
      RECT 10.855 2.34 11.025 3.075 ;
      RECT 8.735 2.265 9.065 3.075 ;
      RECT 10.175 2.34 10.345 3.075 ;
      RECT 11.535 2.34 11.705 3.075 ;
      RECT 7.195 1.425 7.525 2.735 ;
      RECT 10.855 2.34 11.705 2.51 ;
      RECT 8.735 2.34 10.345 2.51 ;
      RECT 7.195 2.265 9.065 2.435 ;
      RECT 8.55 1.425 8.88 1.755 ;
      RECT 7.04 1.425 8.88 1.595 ;
      RECT 7.04 0.595 7.21 1.595 ;
      RECT 6.88 0.595 7.21 0.925 ;
      RECT 11.875 2 12.125 2.575 ;
      RECT 11.52 2 12.125 2.17 ;
      RECT 11.52 0.82 11.69 2.17 ;
      RECT 9.59 0.745 9.92 1.12 ;
      RECT 11.145 0.82 11.69 0.99 ;
      RECT 8.97 0.745 10.475 0.915 ;
      RECT 11.145 0.595 11.315 0.99 ;
      RECT 10.305 0.595 11.315 0.765 ;
      RECT 8.97 0.585 9.3 0.915 ;
      RECT 10.515 2 10.685 2.735 ;
      RECT 9.235 2 11.35 2.17 ;
      RECT 11.18 1.16 11.35 2.17 ;
      RECT 8.01 1.925 9.405 2.095 ;
      RECT 8.01 1.765 8.34 2.095 ;
      RECT 10.645 1.16 11.35 1.33 ;
      RECT 10.645 0.935 10.975 1.33 ;
      RECT 3.205 2.405 3.925 2.735 ;
      RECT 3.205 1.98 3.455 2.735 ;
      RECT 3 1.98 3.455 2.15 ;
      RECT 3 0.255 3.17 2.15 ;
      RECT 9.09 1.085 9.42 1.725 ;
      RECT 5.95 1.095 6.54 1.425 ;
      RECT 7.38 1.085 9.42 1.255 ;
      RECT 5.95 0.255 6.12 1.425 ;
      RECT 7.38 0.255 7.78 1.255 ;
      RECT 4.405 0.615 5.44 0.785 ;
      RECT 5.27 0.255 5.44 0.785 ;
      RECT 2.825 0.255 3.17 0.675 ;
      RECT 4.405 0.255 4.575 0.785 ;
      RECT 2.825 0.255 3.57 0.585 ;
      RECT 5.27 0.255 7.78 0.425 ;
      RECT 2.825 0.255 4.575 0.425 ;
      RECT 5.995 2.905 8.34 3.075 ;
      RECT 8.01 2.745 8.34 3.075 ;
      RECT 4.595 1.725 4.925 3.075 ;
      RECT 5.995 2.625 6.165 3.075 ;
      RECT 4.595 2.625 6.165 2.795 ;
      RECT 3.985 1.725 5.44 1.895 ;
      RECT 5.11 1.295 5.44 1.895 ;
      RECT 3.985 0.675 4.235 1.895 ;
      RECT 6.335 2.105 6.665 2.735 ;
      RECT 5.29 2.105 6.665 2.455 ;
      RECT 5.61 0.595 5.78 2.455 ;
      RECT 4.57 0.955 4.9 1.555 ;
      RECT 4.57 0.955 5.78 1.125 ;
      RECT 2.82 2.905 4.425 3.075 ;
      RECT 4.095 2.065 4.425 3.075 ;
      RECT 1.385 2.32 1.715 3.045 ;
      RECT 2.82 2.32 2.99 3.075 ;
      RECT 1.385 2.32 2.99 2.49 ;
      RECT 2.66 1.01 2.83 2.49 ;
      RECT 3.635 2.065 4.425 2.235 ;
      RECT 3.635 0.755 3.805 2.235 ;
      RECT 2.485 1.01 2.83 1.18 ;
      RECT 3.475 0.755 3.805 1.135 ;
      RECT 2.135 0.84 2.655 1.01 ;
      RECT 2.135 0.5 2.305 1.01 ;
      RECT 1.525 0.5 2.305 0.67 ;
      RECT 1.525 0.255 1.855 0.67 ;
      RECT 0.085 1.91 0.385 3.045 ;
      RECT 0.085 1.91 1.905 2.08 ;
      RECT 0.585 1.75 1.905 2.08 ;
      RECT 0.085 0.255 0.255 3.045 ;
      RECT 0.585 1.555 0.915 2.08 ;
      RECT 0.085 0.255 0.415 0.675 ;
  END
END scs130lp_srsdfxtp_1

MACRO scs130lp_tap_1
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_tap_1 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0.09 0.265 0.39 1.44 ;
    END
  END vnb
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 1.89 0.39 3.065 ;
    END
  END vpb
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.48 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.48 3.415 ;
    END
  END vpwr
END scs130lp_tap_1

MACRO scs130lp_tap_2
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_tap_2 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0.09 0.265 0.87 1.44 ;
    END
  END vnb
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 1.89 0.87 3.065 ;
    END
  END vpb
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
      LAYER li ;
        RECT 0 -0.085 0.96 0.085 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
      LAYER li ;
        RECT 0 3.245 0.96 3.415 ;
    END
  END vpwr
END scs130lp_tap_2

MACRO scs130lp_tapvgnd2_1
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_tapvgnd2_1 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 0.48 0.085 ;
        RECT 0.09 -0.085 0.39 1.44 ;
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 1.89 0.39 3.065 ;
      LAYER met1 ;
        RECT 0.095 2.29 0.385 2.52 ;
    END
  END vpb
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 0.48 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr
END scs130lp_tapvgnd2_1

MACRO scs130lp_tapvgnd_1
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_tapvgnd_1 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 0.48 0.085 ;
        RECT 0.09 -0.085 0.39 1.44 ;
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0.09 1.89 0.39 3.065 ;
      LAYER met1 ;
        RECT 0.095 2.66 0.385 2.89 ;
    END
  END vpb
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 0.48 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr
END scs130lp_tapvgnd_1

MACRO scs130lp_tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_tapvpwrvgnd_1 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li ;
        RECT 0 -0.085 0.48 0.085 ;
        RECT 0.09 -0.085 0.39 1.105 ;
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li ;
        RECT 0 3.245 0.48 3.415 ;
        RECT 0.09 2.205 0.39 3.415 ;
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr
END scs130lp_tapvpwrvgnd_1

MACRO scs130lp_xnor2_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor2_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.545 0.255 1.34 0.515 ;
        RECT 0.545 0.255 0.715 2.095 ;
        RECT 0.085 1.43 0.57 2.245 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.305 1.425 2.455 1.895 ;
        RECT 1.595 1.22 2.455 1.895 ;
        RECT 1.305 1.425 1.57 2.095 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3033 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.27 2.405 3.27 2.575 ;
        RECT 3.1 0.345 3.27 2.575 ;
        RECT 2.75 0.345 3.27 1.38 ;
        RECT 2.27 2.405 2.6 3.025 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.925 -0.085 2.18 0.675 ;
        RECT 0.095 -0.085 0.375 1.26 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.77 2.745 3.06 3.415 ;
        RECT 1.16 2.605 1.79 3.415 ;
        RECT 0.26 2.415 0.57 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.74 2.265 0.99 3.065 ;
      RECT 0.74 2.265 2.1 2.435 ;
      RECT 1.93 2.065 2.1 2.435 ;
      RECT 0.885 0.93 1.125 2.435 ;
      RECT 1.93 2.065 2.93 2.235 ;
      RECT 2.67 1.565 2.93 2.235 ;
      RECT 0.885 0.93 1.215 1.26 ;
      RECT 1.51 0.845 2.58 1.035 ;
      RECT 2.35 0.345 2.58 1.035 ;
      RECT 1.51 0.345 1.755 1.035 ;
  END
END scs130lp_xnor2_0

MACRO scs130lp_xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor2_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.425 1.655 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.825 1.425 2.465 1.845 ;
        RECT 0.085 1.92 1.995 2.09 ;
        RECT 1.825 1.425 1.995 2.09 ;
        RECT 0.085 1.185 0.44 2.09 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6573 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 2.355 3.275 2.555 ;
        RECT 3.095 0.255 3.275 2.555 ;
        RECT 3.015 1.845 3.275 2.555 ;
        RECT 3.015 0.255 3.275 1.175 ;
        RECT 2.505 2.355 2.765 3.075 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.97 -0.085 2.3 0.575 ;
        RECT 0.95 -0.085 1.28 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.935 2.725 3.265 3.415 ;
        RECT 0.985 2.6 1.825 3.415 ;
        RECT 0.125 2.26 0.385 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.555 2.26 0.815 3.075 ;
      RECT 0.555 2.26 2.335 2.43 ;
      RECT 2.165 2.015 2.335 2.43 ;
      RECT 2.165 2.015 2.845 2.185 ;
      RECT 2.675 1.085 2.845 2.185 ;
      RECT 2.675 1.345 2.925 1.675 ;
      RECT 0.61 1.085 2.845 1.255 ;
      RECT 0.61 0.845 0.78 1.255 ;
      RECT 0.125 0.845 0.78 1.015 ;
      RECT 0.125 0.265 0.455 1.015 ;
      RECT 1.47 0.745 2.835 0.915 ;
      RECT 2.505 0.255 2.835 0.915 ;
      RECT 1.47 0.255 1.8 0.915 ;
  END
END scs130lp_xnor2_1

MACRO scs130lp_xnor2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor2_2 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.465 1.405 3.135 1.575 ;
        RECT 2.465 1.005 2.635 1.575 ;
        RECT 1.655 1.005 2.635 1.175 ;
        RECT 1.02 1.425 1.825 1.75 ;
        RECT 1.655 1.005 1.825 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.305 1.405 4.5 1.75 ;
        RECT 2.115 1.745 3.475 1.915 ;
        RECT 2.115 1.345 2.285 1.915 ;
        RECT 1.995 1.345 2.285 1.675 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2558 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.885 1.065 6.155 3.075 ;
        RECT 5.025 1.775 6.155 1.945 ;
        RECT 5.315 1.065 6.155 1.235 ;
        RECT 5.315 0.595 5.645 1.235 ;
        RECT 5.025 1.775 5.215 3.075 ;
        RECT 4.095 2.26 5.215 2.43 ;
        RECT 4.095 2.26 4.355 2.635 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 4.025 -0.085 4.785 0.895 ;
        RECT 3.165 -0.085 3.495 0.895 ;
        RECT 0.585 -0.085 0.805 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.385 2.115 5.715 3.415 ;
        RECT 3.2 2.775 3.46 3.415 ;
        RECT 2.195 2.435 2.525 3.415 ;
        RECT 1.235 2.26 1.565 3.415 ;
        RECT 0.3 2.27 0.645 3.415 ;
        RECT 0.3 1.815 0.51 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.805 1.065 5.145 1.235 ;
      RECT 4.955 0.255 5.145 1.235 ;
      RECT 3.665 0.3 3.855 1.235 ;
      RECT 2.805 0.3 2.995 1.235 ;
      RECT 5.815 0.255 6.145 0.895 ;
      RECT 4.955 0.255 6.145 0.425 ;
      RECT 1.745 2.085 2.015 3.075 ;
      RECT 0.815 1.92 1.065 3.075 ;
      RECT 1.745 2.085 3.855 2.255 ;
      RECT 0.68 1.075 0.85 2.1 ;
      RECT 4.685 1.405 4.855 2.09 ;
      RECT 3.645 1.92 4.855 2.09 ;
      RECT 0.68 1.92 1.945 2.09 ;
      RECT 4.685 1.405 5.715 1.605 ;
      RECT 0.68 1.075 1.485 1.245 ;
      RECT 1.315 0.615 1.485 1.245 ;
      RECT 1.315 0.615 2.015 0.815 ;
      RECT 2.7 2.435 3.03 3.075 ;
      RECT 3.63 2.895 4.855 3.065 ;
      RECT 4.525 2.6 4.855 3.065 ;
      RECT 3.63 2.435 3.855 3.065 ;
      RECT 2.7 2.435 3.855 2.605 ;
      RECT 0.095 0.735 0.425 1.095 ;
      RECT 0.095 0.735 1.145 0.905 ;
      RECT 0.975 0.255 1.145 0.905 ;
      RECT 2.185 0.255 2.515 0.835 ;
      RECT 0.095 0.255 0.415 1.095 ;
      RECT 0.975 0.255 2.515 0.445 ;
  END
END scs130lp_xnor2_2

MACRO scs130lp_xnor2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor2_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.52 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.305 1.425 7.96 1.595 ;
        RECT 6.305 1.425 6.475 1.935 ;
        RECT 3.5 1.765 6.475 1.935 ;
        RECT 3.5 1.415 3.83 1.935 ;
        RECT 1.285 1.93 3.67 2.1 ;
        RECT 1.285 1.415 1.57 2.1 ;
        RECT 0.445 1.415 1.57 1.75 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9404 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.82 2.105 6.08 3.075 ;
        RECT 4.165 2.105 6.08 2.275 ;
        RECT 0.095 1.075 5.435 1.245 ;
        RECT 5.105 0.595 5.435 1.245 ;
        RECT 4.215 2.105 4.645 3.075 ;
        RECT 4.235 0.605 4.435 1.245 ;
        RECT 0.945 2.27 4.645 2.45 ;
        RECT 0.945 1.92 1.115 2.45 ;
        RECT 0.095 1.92 1.115 2.09 ;
        RECT 0.095 1.075 0.275 2.09 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
      ANTENNAGATEAREA 2.52 LAYER met1 ;
      ANTENNAMAXAREACAR 0.348214 LAYER li ;
      ANTENNAMAXAREACAR 0.348214 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.26746 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.26746 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.022937 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 8.255 1.55 8.545 1.78 ;
        RECT 2.015 1.595 8.545 1.735 ;
        RECT 2.015 1.55 2.305 1.78 ;
      LAYER li ;
        RECT 8.24 1.425 9.59 1.75 ;
        RECT 2.075 1.415 3.16 1.75 ;
        RECT 1.81 1.415 3.16 1.595 ;
    END
  END B
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 7.505 -0.085 7.835 0.575 ;
        RECT 6.635 -0.085 6.965 0.575 ;
        RECT 3.225 -0.085 3.555 0.565 ;
        RECT 2.365 -0.085 2.695 0.565 ;
        RECT 1.505 -0.085 1.835 0.565 ;
        RECT 0.635 -0.085 0.965 0.565 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 9.62 2.26 9.95 3.415 ;
        RECT 8.76 2.26 9.09 3.415 ;
        RECT 7.9 2.26 8.23 3.415 ;
        RECT 7.04 2.125 7.37 3.415 ;
        RECT 6.25 2.125 6.47 3.415 ;
        RECT 4.815 2.445 5.65 3.415 ;
        RECT 3.715 2.62 4.045 3.415 ;
        RECT 1.035 2.96 1.365 3.415 ;
        RECT 0.095 2.26 0.425 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 9.26 1.92 9.45 3.075 ;
      RECT 8.4 1.92 8.59 3.075 ;
      RECT 7.54 1.775 7.73 3.075 ;
      RECT 6.645 1.775 6.87 3.075 ;
      RECT 7.54 1.92 9.99 2.09 ;
      RECT 9.77 1.065 9.99 2.09 ;
      RECT 6.645 1.775 7.8 1.945 ;
      RECT 4.04 1.415 6.135 1.585 ;
      RECT 5.625 1.085 6.135 1.585 ;
      RECT 5.625 1.085 9.99 1.255 ;
      RECT 8.365 1.065 9.99 1.255 ;
      RECT 9.225 0.615 9.555 1.255 ;
      RECT 8.365 0.615 8.695 1.255 ;
      RECT 6.135 0.745 8.195 0.915 ;
      RECT 8.005 0.255 8.195 0.915 ;
      RECT 9.725 0.255 9.985 0.895 ;
      RECT 8.865 0.255 9.055 0.895 ;
      RECT 7.135 0.285 7.335 0.915 ;
      RECT 6.135 0.305 6.465 0.915 ;
      RECT 8.005 0.255 9.055 0.435 ;
      RECT 8.005 0.255 9.985 0.425 ;
      RECT 5.605 0.255 5.935 0.915 ;
      RECT 4.605 0.255 4.935 0.905 ;
      RECT 0.135 0.735 4.065 0.905 ;
      RECT 3.735 0.255 4.065 0.905 ;
      RECT 2.865 0.285 3.055 0.905 ;
      RECT 2.005 0.285 2.195 0.905 ;
      RECT 1.155 0.285 1.335 0.905 ;
      RECT 0.135 0.295 0.465 0.905 ;
      RECT 3.735 0.255 4.935 0.435 ;
      RECT 3.735 0.255 5.935 0.425 ;
      RECT 1.535 2.62 3.545 2.96 ;
      RECT 0.595 2.62 0.865 2.95 ;
      RECT 0.595 2.62 3.545 2.79 ;
  END
END scs130lp_xnor2_4

MACRO scs130lp_xnor2_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor2_lp 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.015 1.245 2.345 1.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.626 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.525 1.51 2.92 1.84 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3955 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.845 1.975 1.175 3.065 ;
        RECT 0.105 1.975 1.175 2.145 ;
        RECT 0.105 0.44 0.435 0.9 ;
        RECT 0.105 0.44 0.355 2.145 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.095 -0.085 2.345 1.065 ;
        RECT 1.075 -0.085 1.405 0.935 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.925 2.37 3.255 3.415 ;
        RECT 1.865 2.37 2.195 3.415 ;
        RECT 0.315 2.325 0.645 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.395 2.02 2.725 3.065 ;
      RECT 1.355 2.02 3.27 2.19 ;
      RECT 3.1 0.605 3.27 2.19 ;
      RECT 1.355 1.465 1.525 2.19 ;
      RECT 0.54 1.465 1.525 1.795 ;
      RECT 2.915 0.605 3.27 1.065 ;
      RECT 0.615 1.115 1.835 1.285 ;
      RECT 1.585 0.605 1.835 1.285 ;
      RECT 0.615 0.44 0.865 1.285 ;
  END
END scs130lp_xnor2_lp

MACRO scs130lp_xnor2_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor2_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.21 1.765 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 2.69 2.725 2.97 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4263 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.49 0.62 2.82 0.83 ;
        RECT 2.225 2.28 2.725 2.49 ;
        RECT 2.555 0.62 2.725 2.49 ;
    END
  END Y
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 1.09 0.86 2.3 1.03 ;
        RECT 1.97 0.62 2.3 1.03 ;
        RECT 1.09 -0.085 1.28 1.03 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 2.905 2.18 3.095 3.415 ;
        RECT 1.1 2.28 1.43 2.49 ;
        RECT 1.1 2.28 1.27 3.415 ;
        RECT 0.24 2.28 0.57 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 3 0.27 3.19 0.76 ;
      RECT 1.46 0.27 1.79 0.68 ;
      RECT 1.46 0.27 3.19 0.44 ;
      RECT 0.75 1.93 0.92 2.42 ;
      RECT 0.24 1.93 2.375 2.1 ;
      RECT 2.205 1.28 2.375 2.1 ;
      RECT 0.24 0.62 0.41 2.1 ;
      RECT 0.24 0.62 0.57 0.83 ;
  END
END scs130lp_xnor2_m

MACRO scs130lp_xnor3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor3_1 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.246 LAYER li ;
    PORT
      LAYER li ;
        RECT 6.845 1.18 7.185 1.51 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.729 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.515 1.345 3.845 1.78 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.381 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.025 1.345 1.315 1.78 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5754 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.1 0.255 0.44 1.125 ;
        RECT 0.1 1.815 0.35 3.075 ;
        RECT 0.1 0.255 0.27 3.075 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
      LAYER li ;
        RECT 0 -0.085 8.16 0.085 ;
        RECT 7.115 -0.085 7.445 0.605 ;
        RECT 3.305 -0.085 3.635 0.445 ;
        RECT 0.65 -0.085 0.98 0.365 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
      LAYER li ;
        RECT 0 3.245 8.16 3.415 ;
        RECT 7.16 2.345 7.49 3.415 ;
        RECT 3.315 2.865 3.645 3.415 ;
        RECT 0.53 2.29 0.78 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 7.775 2.29 8.065 2.52 ;
      RECT 5.375 2.29 5.665 2.52 ;
      RECT 5.375 2.335 8.065 2.475 ;
      RECT 4.895 1.18 5.185 1.41 ;
      RECT 2.495 1.18 2.785 1.41 ;
      RECT 2.495 1.225 5.185 1.365 ;
    LAYER li ;
      RECT 7.695 1.895 8.075 2.935 ;
      RECT 7.835 0.34 8.075 2.935 ;
      RECT 7.695 0.34 8.075 1.02 ;
      RECT 4.335 2.895 6.945 3.065 ;
      RECT 6.615 1.845 6.945 3.065 ;
      RECT 4.335 2.71 4.665 3.065 ;
      RECT 6.615 1.845 7.525 2.175 ;
      RECT 7.355 0.775 7.525 2.175 ;
      RECT 7.355 1.19 7.645 1.52 ;
      RECT 6.615 0.775 7.525 0.945 ;
      RECT 6.615 0.255 6.945 0.945 ;
      RECT 4.41 0.255 4.74 0.445 ;
      RECT 4.41 0.255 6.945 0.425 ;
      RECT 5.425 2.515 6.445 2.685 ;
      RECT 6.275 1.115 6.445 2.685 ;
      RECT 5.425 1.845 5.755 2.685 ;
      RECT 6.275 1.115 6.565 1.675 ;
      RECT 5.455 1.115 6.565 1.285 ;
      RECT 5.455 0.935 5.785 1.285 ;
      RECT 4.88 1.875 5.21 2.725 ;
      RECT 1.825 2.525 3.345 2.695 ;
      RECT 3.175 0.615 3.345 2.695 ;
      RECT 3.175 2.37 5.21 2.54 ;
      RECT 1.825 2.235 2.075 2.695 ;
      RECT 2.745 0.615 3.345 1.01 ;
      RECT 6.115 0.595 6.445 0.94 ;
      RECT 2.745 0.615 5.08 0.785 ;
      RECT 4.91 0.595 6.445 0.765 ;
      RECT 2.745 0.525 3.075 1.01 ;
      RECT 5.935 1.455 6.105 2.345 ;
      RECT 4.955 1.455 6.105 1.625 ;
      RECT 4.955 0.955 5.285 1.625 ;
      RECT 4.925 0.955 5.285 1.205 ;
      RECT 3.745 2.03 4.66 2.2 ;
      RECT 4.49 1.375 4.66 2.2 ;
      RECT 3.745 1.95 4.185 2.2 ;
      RECT 4.015 0.955 4.185 2.2 ;
      RECT 4.49 1.375 4.785 1.705 ;
      RECT 3.85 0.955 4.185 1.125 ;
      RECT 2.835 1.18 3.005 2.355 ;
      RECT 1.825 1.18 3.005 1.385 ;
      RECT 1.825 0.875 2.075 1.385 ;
      RECT 1.29 1.95 1.655 2.495 ;
      RECT 1.485 0.875 1.655 2.495 ;
      RECT 1.485 1.555 2.665 1.885 ;
      RECT 1.195 0.875 1.655 1.125 ;
      RECT 0.95 2.865 2.505 3.035 ;
      RECT 0.95 1.95 1.12 3.035 ;
      RECT 0.61 1.95 1.12 2.12 ;
      RECT 0.61 0.535 0.78 2.12 ;
      RECT 0.44 1.295 0.78 1.625 ;
      RECT 2.245 0.525 2.575 1.01 ;
      RECT 0.61 0.535 2.575 0.705 ;
  END
END scs130lp_xnor3_1

MACRO scs130lp_xnor3_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xnor3_lp 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.465 1.515 0.835 1.845 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.002 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.045 1.345 3.03 1.78 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.73 0.975 8.06 1.38 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.375 1.18 9.965 2.89 ;
        RECT 9.715 0.64 9.965 2.89 ;
        RECT 9.375 1.18 9.705 3.025 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 8.845 0.73 9.535 0.9 ;
        RECT 9.365 -0.085 9.535 0.9 ;
        RECT 8.845 0.73 9.175 1.1 ;
        RECT 2.475 -0.085 2.725 0.815 ;
        RECT 0.905 -0.085 1.155 0.985 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 8.845 1.985 9.175 3.415 ;
        RECT 2.6 2.595 2.93 3.415 ;
        RECT 0.77 2.025 1.1 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 6.715 1.645 7.185 1.975 ;
      RECT 6.715 0.265 6.965 1.975 ;
      RECT 8.855 0.265 9.185 0.55 ;
      RECT 6.715 0.265 9.185 0.435 ;
      RECT 8.315 1.56 8.645 3.025 ;
      RECT 8.475 0.615 8.645 3.025 ;
      RECT 8.05 1.56 8.645 1.795 ;
      RECT 7.715 0.615 8.645 0.795 ;
      RECT 3.795 2.895 8.065 3.065 ;
      RECT 7.895 1.975 8.065 3.065 ;
      RECT 6.325 2.505 6.655 3.065 ;
      RECT 4.915 1.795 5.085 3.065 ;
      RECT 3.795 2.595 4.125 3.065 ;
      RECT 7.365 1.975 8.065 2.145 ;
      RECT 7.365 0.615 7.535 2.145 ;
      RECT 4.915 1.795 5.615 1.965 ;
      RECT 5.285 0.965 5.615 1.965 ;
      RECT 7.145 0.615 7.535 0.995 ;
      RECT 5.265 2.145 5.595 2.715 ;
      RECT 7.465 2.325 7.715 2.685 ;
      RECT 6.835 2.325 7.715 2.495 ;
      RECT 5.265 2.155 7.005 2.325 ;
      RECT 6.305 0.265 6.475 2.325 ;
      RECT 4.075 0.265 4.245 0.715 ;
      RECT 4.075 0.265 6.475 0.435 ;
      RECT 0.115 2.025 0.57 3.065 ;
      RECT 0.115 0.525 0.285 3.065 ;
      RECT 5.795 0.615 6.125 1.965 ;
      RECT 1.175 1.165 1.505 1.835 ;
      RECT 1.335 0.265 1.505 1.835 ;
      RECT 0.115 1.165 1.505 1.335 ;
      RECT 2.125 0.995 3.075 1.165 ;
      RECT 2.905 0.265 3.075 1.165 ;
      RECT 0.115 0.525 0.445 1.335 ;
      RECT 3.725 0.895 4.595 1.065 ;
      RECT 4.425 0.615 4.595 1.065 ;
      RECT 2.125 0.265 2.295 1.165 ;
      RECT 3.725 0.265 3.895 1.065 ;
      RECT 4.425 0.615 6.125 0.785 ;
      RECT 2.905 0.265 3.895 0.435 ;
      RECT 1.335 0.265 2.295 0.435 ;
      RECT 1.3 2.025 1.63 3.065 ;
      RECT 4.405 1.245 4.735 2.715 ;
      RECT 1.3 2.245 4.735 2.415 ;
      RECT 1.3 2.025 1.865 2.415 ;
      RECT 1.695 0.615 1.865 2.415 ;
      RECT 4.405 1.245 5.105 1.415 ;
      RECT 4.775 0.965 5.105 1.415 ;
      RECT 1.695 0.615 1.945 0.985 ;
      RECT 3.21 1.815 3.54 2.065 ;
      RECT 3.295 0.615 3.54 2.065 ;
      RECT 3.295 1.245 3.83 1.575 ;
      RECT 3.295 0.615 3.545 1.575 ;
  END
END scs130lp_xnor3_lp

MACRO scs130lp_xor2_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor2_0 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.21 1.35 1.395 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.205 1.565 1.94 1.855 ;
        RECT 1.52 1.21 1.94 1.855 ;
        RECT 0.205 1.185 0.455 1.855 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5161 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.545 1.815 2.815 2.495 ;
        RECT 2.645 0.41 2.815 2.495 ;
        RECT 1.97 0.41 2.815 0.7 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.985 -0.085 3.255 0.8 ;
        RECT 1.13 -0.085 1.46 0.7 ;
        RECT 0.27 -0.085 0.56 0.8 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.81 2.705 2.035 3.415 ;
        RECT 0.915 2.385 1.21 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.38 2.365 1.64 3.065 ;
      RECT 2.205 2.665 3.255 2.835 ;
      RECT 2.985 1.815 3.255 2.835 ;
      RECT 2.205 2.365 2.375 2.835 ;
      RECT 1.38 2.365 2.375 2.535 ;
      RECT 0.095 2.025 0.425 3.065 ;
      RECT 0.095 2.025 2.375 2.195 ;
      RECT 2.205 0.87 2.375 2.195 ;
      RECT 2.205 0.87 2.475 1.625 ;
      RECT 0.73 0.87 2.475 1.04 ;
      RECT 0.73 0.395 0.96 1.04 ;
  END
END scs130lp_xor2_0

MACRO scs130lp_xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor2_1 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.625 1.21 1.765 1.555 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.085 1.725 2.115 1.895 ;
        RECT 1.935 1.345 2.115 1.895 ;
        RECT 0.085 1.21 0.455 1.895 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8463 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.505 1.795 2.835 2.065 ;
        RECT 2.505 1.57 2.735 2.065 ;
        RECT 2.285 1.57 2.735 1.75 ;
        RECT 2.285 0.595 2.455 1.75 ;
        RECT 2.04 0.595 2.455 1.165 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.965 -0.085 3.215 1.06 ;
        RECT 1.03 -0.085 1.36 0.7 ;
        RECT 0.17 -0.085 0.43 1.04 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.965 2.915 2.295 3.415 ;
        RECT 0.99 2.405 1.27 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 1.44 2.405 1.77 3.075 ;
      RECT 2.935 2.575 3.265 2.925 ;
      RECT 1.44 2.575 3.265 2.745 ;
      RECT 0.17 2.065 0.5 3.075 ;
      RECT 1.94 2.235 3.235 2.405 ;
      RECT 3.065 1.23 3.235 2.405 ;
      RECT 0.17 2.065 2.11 2.235 ;
      RECT 2.905 1.23 3.235 1.625 ;
      RECT 2.625 1.23 3.235 1.4 ;
      RECT 2.625 0.255 2.795 1.4 ;
      RECT 0.6 0.87 1.87 1.04 ;
      RECT 1.7 0.255 1.87 1.04 ;
      RECT 0.6 0.335 0.86 1.04 ;
      RECT 1.7 0.255 2.795 0.425 ;
  END
END scs130lp_xor2_1

MACRO scs130lp_xor2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor2_2 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.9 1.92 5.725 2.09 ;
        RECT 5.395 1.415 5.725 2.09 ;
        RECT 3.9 1.355 4.07 2.09 ;
        RECT 3.74 0.615 3.92 1.605 ;
        RECT 0.37 0.615 3.92 0.785 ;
        RECT 0.675 1.95 2.335 2.12 ;
        RECT 1.595 1.345 2.335 2.12 ;
        RECT 0.675 1.345 0.845 2.12 ;
        RECT 0.37 1.345 0.845 1.605 ;
        RECT 0.37 0.615 0.54 1.605 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8442 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.05 2.26 6.155 2.43 ;
        RECT 5.895 1.075 6.155 2.43 ;
        RECT 4.475 1.075 6.155 1.245 ;
        RECT 4.475 0.81 5.125 1.245 ;
        RECT 4.475 0.595 4.805 1.245 ;
        RECT 3.05 1.84 3.38 2.43 ;
        RECT 3.21 0.955 3.38 2.43 ;
        RECT 3.025 0.955 3.38 1.16 ;
    END
  END X
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.63 LAYER li ;
      ANTENNAGATEAREA 1.26 LAYER met1 ;
      ANTENNAMAXAREACAR 0.35627 LAYER li ;
      ANTENNAMAXAREACAR 0.35627 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.319048 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.319048 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.045873 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 4.415 1.55 4.705 1.78 ;
        RECT 1.055 1.595 4.705 1.735 ;
        RECT 1.055 1.55 1.345 1.78 ;
      LAYER li ;
        RECT 4.285 1.415 4.955 1.75 ;
        RECT 1.015 1.345 1.425 1.78 ;
    END
  END B
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
      LAYER li ;
        RECT 0 -0.085 6.24 0.085 ;
        RECT 5.795 -0.085 6.125 0.905 ;
        RECT 3.535 -0.085 3.865 0.445 ;
        RECT 2.48 -0.085 2.81 0.445 ;
        RECT 1.23 -0.085 1.56 0.445 ;
        RECT 0.195 -0.085 0.525 0.445 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
      LAYER li ;
        RECT 0 3.245 6.24 3.415 ;
        RECT 5.01 2.94 5.34 3.415 ;
        RECT 3.99 2.94 4.32 3.415 ;
        RECT 2.1 2.63 2.43 3.415 ;
        RECT 0.255 2.29 0.62 3.415 ;
        RECT 0.255 1.82 0.505 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.62 2.63 3.81 3.075 ;
      RECT 2.965 2.6 5.85 2.77 ;
      RECT 4.09 0.255 4.305 1.185 ;
      RECT 5.295 0.255 5.625 0.905 ;
      RECT 4.975 0.255 5.625 0.64 ;
      RECT 4.09 0.255 5.625 0.425 ;
      RECT 1.19 2.29 1.43 2.63 ;
      RECT 1.19 2.29 2.7 2.46 ;
      RECT 2.53 0.955 2.7 2.46 ;
      RECT 2.53 1.33 3.03 1.605 ;
      RECT 0.72 0.955 2.7 1.175 ;
      RECT 0.79 2.8 1.93 3.075 ;
      RECT 1.6 2.63 1.93 3.075 ;
      RECT 0.79 2.29 1.02 3.075 ;
  END
END scs130lp_xor2_2

MACRO scs130lp_xor2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor2_4 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6464 LAYER li ;
    PORT
      LAYER li ;
        RECT 3.995 2.29 5.195 2.605 ;
        RECT 4.865 1.845 5.195 2.605 ;
        RECT 3.995 1.015 5.155 1.185 ;
        RECT 4.965 0.255 5.155 1.185 ;
        RECT 4.105 0.255 4.295 1.185 ;
        RECT 3.995 0.695 4.275 2.605 ;
        RECT 1.815 0.695 4.295 0.905 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
      ANTENNAGATEAREA 2.52 LAYER met1 ;
      ANTENNAMAXAREACAR 0.615397 LAYER li ;
      ANTENNAMAXAREACAR 0.615397 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.623016 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.623016 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.045873 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 6.335 1.18 6.625 1.41 ;
        RECT 1.26 1.225 6.625 1.365 ;
        RECT 3.455 1.18 3.745 1.41 ;
        RECT 1.26 1.18 1.55 1.41 ;
      LAYER li ;
        RECT 6.305 1.355 7.655 1.535 ;
        RECT 6.305 1.2 7.075 1.535 ;
        RECT 3.34 1.075 3.685 1.435 ;
        RECT 1.26 1.075 3.685 1.245 ;
        RECT 0.4 1.275 1.555 1.525 ;
        RECT 1.26 1.075 1.555 1.525 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.26 LAYER li ;
      ANTENNAGATEAREA 2.52 LAYER met1 ;
      ANTENNAMAXAREACAR 0.385714 LAYER li ;
      ANTENNAMAXAREACAR 0.385714 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.352381 LAYER li ;
      ANTENNAMAXSIDEAREACAR 0.352381 LAYER met1 ;
      ANTENNAMAXCUTCAR 0.022937 LAYER mcon ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.55 8.065 1.78 ;
        RECT 2.495 1.595 8.065 1.735 ;
        RECT 2.495 1.55 2.785 1.78 ;
      LAYER li ;
        RECT 7.825 1.355 9.6 1.535 ;
        RECT 7.825 1.355 8.015 1.8 ;
        RECT 1.735 1.415 3.085 1.775 ;
    END
  END B
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
      LAYER li ;
        RECT 0 -0.085 10.08 0.085 ;
        RECT 9.325 -0.085 9.655 0.845 ;
        RECT 8.465 -0.085 8.795 0.845 ;
        RECT 7.605 -0.085 7.935 0.845 ;
        RECT 6.745 -0.085 7.075 0.69 ;
        RECT 5.325 -0.085 6.215 0.69 ;
        RECT 5.325 -0.085 5.655 1.105 ;
        RECT 4.465 -0.085 4.795 0.845 ;
        RECT 3.605 -0.085 3.935 0.525 ;
        RECT 0.985 -0.085 1.215 0.565 ;
        RECT 0.095 -0.085 0.425 1.095 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
      LAYER li ;
        RECT 0 3.245 10.08 3.415 ;
        RECT 7.245 2.31 7.575 3.415 ;
        RECT 6.385 2.31 6.715 3.415 ;
        RECT 3.12 2.285 3.45 3.415 ;
        RECT 2.245 2.285 2.575 3.415 ;
        RECT 1.385 2.285 1.715 3.415 ;
        RECT 0.525 2.035 0.855 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 8.965 1.705 9.295 2.735 ;
      RECT 8.185 1.705 8.435 2.735 ;
      RECT 8.185 1.705 9.995 1.875 ;
      RECT 9.77 1.015 9.995 1.875 ;
      RECT 4.445 1.355 6.135 1.535 ;
      RECT 5.825 0.86 6.135 1.535 ;
      RECT 7.245 1.015 9.995 1.185 ;
      RECT 5.825 0.86 7.435 1.03 ;
      RECT 8.965 0.255 9.155 1.185 ;
      RECT 8.105 0.255 8.295 1.185 ;
      RECT 7.245 0.255 7.435 1.185 ;
      RECT 6.385 0.255 6.575 1.03 ;
      RECT 7.745 2.905 9.725 3.075 ;
      RECT 9.465 2.045 9.725 3.075 ;
      RECT 6.885 1.97 7.075 3.075 ;
      RECT 5.955 1.97 6.215 3.075 ;
      RECT 8.605 2.045 8.795 3.075 ;
      RECT 7.745 1.97 7.935 3.075 ;
      RECT 5.955 1.97 7.935 2.14 ;
      RECT 3.625 2.775 5.625 3.075 ;
      RECT 5.365 1.815 5.625 3.075 ;
      RECT 2.745 1.945 2.95 3.075 ;
      RECT 1.885 1.945 2.075 3.075 ;
      RECT 1.025 1.695 1.215 3.075 ;
      RECT 0.095 1.695 0.355 3.075 ;
      RECT 3.625 1.945 3.825 3.075 ;
      RECT 1.025 1.945 3.825 2.115 ;
      RECT 1.025 1.695 1.225 2.115 ;
      RECT 0.095 1.695 1.225 1.865 ;
      RECT 0.595 0.255 0.785 1.095 ;
      RECT 0.595 0.735 1.645 0.905 ;
      RECT 1.385 0.255 1.645 0.905 ;
      RECT 0.595 0.255 0.815 0.905 ;
      RECT 1.385 0.255 3.435 0.525 ;
  END
END scs130lp_xor2_4

MACRO scs130lp_xor2_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor2_lp 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.085 1.69 3.265 1.86 ;
        RECT 2.935 1.18 3.265 1.86 ;
        RECT 1.085 1.295 1.9 1.86 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.29 1.18 2.755 1.51 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4176 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.735 0.575 1.235 1.035 ;
        RECT 0.125 1.215 0.905 1.385 ;
        RECT 0.735 0.575 0.905 1.385 ;
        RECT 0.125 2.075 0.555 3.065 ;
        RECT 0.125 1.215 0.355 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.84 0.085 ;
        RECT 3.385 -0.085 3.715 0.65 ;
        RECT 1.775 -0.085 2.105 0.78 ;
        RECT 0.115 -0.085 0.445 1.035 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.84 3.415 ;
        RECT 3.385 2.39 3.715 3.415 ;
        RECT 1.3 2.74 1.63 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 2.395 2.04 2.725 3.065 ;
      RECT 0.735 2.04 3.615 2.21 ;
      RECT 3.445 0.83 3.615 2.21 ;
      RECT 0.735 1.565 0.905 2.21 ;
      RECT 0.535 1.565 0.905 1.895 ;
      RECT 2.595 0.83 3.615 1 ;
      RECT 2.595 0.32 2.925 1 ;
      RECT 1.83 2.39 2.16 3.065 ;
      RECT 0.77 2.39 1.1 3.065 ;
      RECT 0.77 2.39 2.16 2.56 ;
  END
END scs130lp_xor2_lp

MACRO scs130lp_xor2_m
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor2_m 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.635 1.91 1.285 2.49 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER li ;
    PORT
      LAYER li ;
        RECT 1.595 0.265 2.245 1.38 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3234 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.765 2.625 3.205 2.86 ;
        RECT 3.035 1.21 3.205 2.86 ;
        RECT 2.425 1.21 3.205 1.38 ;
        RECT 2.425 0.89 2.615 1.38 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
      LAYER li ;
        RECT 0 -0.085 3.36 0.085 ;
        RECT 2.87 -0.085 3.2 1.03 ;
        RECT 1.045 -0.085 1.375 1.03 ;
        RECT 0.225 -0.085 0.415 1.09 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
      LAYER li ;
        RECT 0 3.245 3.36 3.415 ;
        RECT 1.875 2.785 2.085 3.415 ;
        RECT 0.955 2.845 1.285 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER li ;
      RECT 0.225 1.56 0.435 3 ;
      RECT 2.685 1.56 2.855 2.23 ;
      RECT 0.225 1.56 2.855 1.73 ;
      RECT 0.655 0.89 0.865 1.73 ;
      RECT 1.465 2.435 1.655 2.985 ;
      RECT 2.335 2.435 2.585 2.765 ;
      RECT 1.465 2.435 2.585 2.605 ;
  END
END scs130lp_xor2_m

MACRO scs130lp_xor3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor3_1 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.246 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.97 1.18 1.3 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.729 LAYER li ;
    PORT
      LAYER li ;
        RECT 5.26 1.18 5.635 1.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.381 LAYER li ;
    PORT
      LAYER li ;
        RECT 7.22 1.18 7.535 1.715 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5985 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.19 0.265 9.475 3.065 ;
        RECT 9.04 0.265 9.475 1.125 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
      LAYER li ;
        RECT 0 -0.085 9.6 0.085 ;
        RECT 8.53 -0.085 8.86 1.125 ;
        RECT 5.61 -0.085 5.86 0.595 ;
        RECT 0.785 -0.085 1.115 0.385 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
      LAYER li ;
        RECT 0 3.245 9.6 3.415 ;
        RECT 8.44 1.815 8.61 3.415 ;
        RECT 5.26 1.765 5.59 3.415 ;
        RECT 0.62 2.195 0.95 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 8.735 1.92 9.025 2.15 ;
      RECT 6.815 1.92 7.105 2.15 ;
      RECT 6.815 1.965 9.025 2.105 ;
      RECT 5.855 1.92 6.145 2.15 ;
      RECT 2.975 1.92 3.265 2.15 ;
      RECT 2.975 1.965 6.145 2.105 ;
    LAYER li ;
      RECT 8.79 1.305 9.01 2.15 ;
      RECT 8.68 1.305 9.01 1.635 ;
      RECT 6.315 2.895 8.235 3.065 ;
      RECT 8.065 0.665 8.235 3.065 ;
      RECT 7.895 2.245 8.235 3.065 ;
      RECT 6.315 1.475 6.645 3.065 ;
      RECT 8.065 0.665 8.315 1.125 ;
      RECT 7.335 1.895 7.715 2.715 ;
      RECT 1.985 2.545 3.71 2.715 ;
      RECT 3.54 0.265 3.71 2.715 ;
      RECT 1.985 2.035 2.315 2.715 ;
      RECT 7.715 0.265 7.885 2.065 ;
      RECT 5.26 0.775 6.34 0.945 ;
      RECT 6.09 0.265 6.34 0.945 ;
      RECT 5.26 0.265 5.43 0.945 ;
      RECT 6.09 0.265 7.885 0.435 ;
      RECT 3.54 0.265 5.43 0.435 ;
      RECT 5.885 1.125 6.135 2.825 ;
      RECT 5.885 1.125 6.69 1.295 ;
      RECT 6.52 0.615 6.69 1.295 ;
      RECT 7.22 0.615 7.47 1 ;
      RECT 6.52 0.615 7.47 0.785 ;
      RECT 6.825 1.92 7.155 2.715 ;
      RECT 6.87 0.965 7.04 2.715 ;
      RECT 4.83 0.615 5.08 3.065 ;
      RECT 3.89 1.395 4.16 1.725 ;
      RECT 3.89 0.615 4.06 1.725 ;
      RECT 3.89 0.615 5.08 0.785 ;
      RECT 1.44 2.895 4.06 3.065 ;
      RECT 3.89 1.905 4.06 3.065 ;
      RECT 1.44 2.015 1.77 3.065 ;
      RECT 3.89 1.905 4.57 2.745 ;
      RECT 4.4 0.965 4.57 2.745 ;
      RECT 0.62 1.845 1.65 2.015 ;
      RECT 0.44 1.525 0.79 1.855 ;
      RECT 1.48 0.915 1.65 3.065 ;
      RECT 4.24 0.965 4.57 1.215 ;
      RECT 3.005 1.865 3.36 2.365 ;
      RECT 3.19 0.265 3.36 2.365 ;
      RECT 2.18 0.265 2.43 1.245 ;
      RECT 2.18 0.265 3.36 0.435 ;
      RECT 0.09 2.035 0.44 3.065 ;
      RECT 2.495 1.425 2.825 2.365 ;
      RECT 2.655 0.615 2.825 2.365 ;
      RECT 0.09 0.565 0.26 3.065 ;
      RECT 1.83 1.425 2.825 1.595 ;
      RECT 1.83 0.565 2 1.595 ;
      RECT 2.655 0.615 3.01 1.245 ;
      RECT 0.09 0.565 0.605 1.245 ;
      RECT 0.09 0.565 2 0.735 ;
  END
END scs130lp_xor3_1

MACRO scs130lp_xor3_lp
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130lp_xor3_lp 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.376 LAYER li ;
    PORT
      LAYER li ;
        RECT 0.835 1.605 1.315 2.15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.002 LAYER li ;
    PORT
      LAYER li ;
        RECT 2.775 1.565 4.425 1.895 ;
        RECT 3.615 1.155 3.945 1.895 ;
        RECT 2.775 1.55 3.235 1.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.689 LAYER li ;
    PORT
      LAYER li ;
        RECT 9.245 1.18 9.955 1.565 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4047 LAYER li ;
    PORT
      LAYER li ;
        RECT 10.675 0.685 10.925 2.89 ;
        RECT 10.125 2.095 10.925 2.265 ;
        RECT 10.125 2.095 10.455 3.065 ;
    END
  END X
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
      LAYER li ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 9.775 0.775 10.495 1 ;
        RECT 10.325 -0.085 10.495 1 ;
        RECT 6.56 -0.085 6.89 0.885 ;
        RECT 1.055 -0.085 1.385 0.915 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
      LAYER li ;
        RECT 0 3.245 11.04 3.415 ;
        RECT 9.595 2.095 9.925 3.415 ;
        RECT 6.26 1.96 6.43 3.415 ;
        RECT 0.855 2.68 1.185 3.415 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
  END vpb
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
  END vnb
  OBS
    LAYER met1 ;
      RECT 7.775 2.29 8.065 2.52 ;
      RECT 4.415 2.29 4.705 2.52 ;
      RECT 4.415 2.335 8.065 2.475 ;
      RECT 4.895 0.81 5.185 1.04 ;
      RECT 2.015 0.81 2.305 1.04 ;
      RECT 2.015 0.855 5.185 0.995 ;
    LAYER li ;
      RECT 7.27 2.895 9.415 3.065 ;
      RECT 9.245 1.745 9.415 3.065 ;
      RECT 7.27 2.01 7.6 3.065 ;
      RECT 9.245 1.745 10.465 1.915 ;
      RECT 10.135 1.235 10.465 1.915 ;
      RECT 7.63 0.265 7.96 1.055 ;
      RECT 9.87 0.265 10.145 0.595 ;
      RECT 7.63 0.265 10.145 0.435 ;
      RECT 7.8 2.01 8.485 2.715 ;
      RECT 8.315 0.615 8.485 2.715 ;
      RECT 8.14 0.615 8.485 1.055 ;
      RECT 6.965 1.5 7.64 1.83 ;
      RECT 7.47 1.235 8.135 1.565 ;
      RECT 4.02 2.895 6.08 3.065 ;
      RECT 5.91 1.15 6.08 3.065 ;
      RECT 6.615 2.01 7.07 3.05 ;
      RECT 4.02 2.075 4.19 3.065 ;
      RECT 2.425 2.075 2.775 2.715 ;
      RECT 2.425 2.075 4.19 2.245 ;
      RECT 2.425 1.185 2.595 2.715 ;
      RECT 6.615 1.15 6.785 3.05 ;
      RECT 2.425 1.185 3.435 1.355 ;
      RECT 3.105 0.615 3.435 1.355 ;
      RECT 5.91 1.15 7.29 1.32 ;
      RECT 7.12 0.595 7.29 1.32 ;
      RECT 7.12 0.595 7.45 1.055 ;
      RECT 5.48 1.45 5.73 2.715 ;
      RECT 5.56 0.265 5.73 2.715 ;
      RECT 5.305 1.45 5.73 1.78 ;
      RECT 5.56 0.425 6.1 0.885 ;
      RECT 5.35 0.265 5.73 0.595 ;
      RECT 4.955 1.96 5.25 2.715 ;
      RECT 4.955 0.575 5.125 2.715 ;
      RECT 4.955 0.575 5.17 1.04 ;
      RECT 4.84 0.575 5.17 1.035 ;
      RECT 4.39 2.31 4.775 2.715 ;
      RECT 4.605 1.215 4.775 2.715 ;
      RECT 4.33 1.215 4.775 1.385 ;
      RECT 4.33 0.31 4.5 1.385 ;
      RECT 4.33 0.31 4.66 1.035 ;
      RECT 1.365 2.895 3.84 3.065 ;
      RECT 3.51 2.425 3.84 3.065 ;
      RECT 0.265 1.095 0.655 3.065 ;
      RECT 1.365 2.33 1.535 3.065 ;
      RECT 0.265 2.33 1.535 2.5 ;
      RECT 0.265 1.095 1.735 1.425 ;
      RECT 1.565 0.265 1.735 1.425 ;
      RECT 0.265 0.545 0.595 3.065 ;
      RECT 3.82 0.265 4.15 0.685 ;
      RECT 1.565 0.265 4.15 0.435 ;
      RECT 1.915 0.81 2.245 2.715 ;
      RECT 1.915 0.81 2.845 1.005 ;
      RECT 2.515 0.625 2.845 1.005 ;
      RECT 8.665 0.685 9.065 2.715 ;
  END
END scs130lp_xor3_lp

END LIBRARY
